-- VHDL produced by vc2vhdl from virtual circuit (vc) description 
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library GhdlLink;
use GhdlLink.LogUtilities.all;
library work;
use work.ahir_system_global_package.all;
entity Inv_Sbox_1_Volatile is -- 
  port ( -- 
    clk, reset: in std_logic; 
    s_in : in  std_logic_vector(7 downto 0);
    s_out : out  std_logic_vector(7 downto 0)-- 
  );
  -- 
end entity Inv_Sbox_1_Volatile;
architecture Inv_Sbox_1_Volatile_arch of Inv_Sbox_1_Volatile is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector(8-1 downto 0);
  signal default_zero_sig: std_logic;
  -- input port buffer signals
  signal s_in_buffer :  std_logic_vector(7 downto 0);
  -- output port buffer signals
  signal s_out_buffer :  std_logic_vector(7 downto 0);
  -- volatile/operator module components. 
  signal global_clock_cycle_count: integer := 0;
  -- 
begin --  
  ---------------------------------------------------------- 
  process(clk)  
  begin -- 
    if(clk'event and clk = '1') then -- 
      if(reset = '1') then -- 
        global_clock_cycle_count <= 0; --
      else -- 
        global_clock_cycle_count <= global_clock_cycle_count + 1; -- 
      end if; --
    end if; --
  end process;
  ---------------------------------------------------------- 
  -- input handling ------------------------------------------------
  s_in_buffer <= s_in;
  -- output handling  -------------------------------------------------------
  s_out <= s_out_buffer;
  -- the control path --------------------------------------------------
  default_zero_sig <= '0';
  -- volatile module, no control path
  -- the data path
  data_path: Block -- 
    signal BITSEL_u8_u1_1004_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1014_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1024_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1034_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1044_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_104_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1054_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1064_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1074_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1084_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1094_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1104_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1114_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1124_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1134_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1144_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_114_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1154_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1164_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1174_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1184_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1194_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1204_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1214_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1224_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1234_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1244_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_124_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1254_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1264_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1274_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1284_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1294_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1302_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1310_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1318_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1326_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1334_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1342_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_134_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1350_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1358_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1366_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1374_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1382_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1390_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1398_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_13_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1406_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1414_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1422_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1430_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1438_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1446_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_144_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1454_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1462_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1470_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1478_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1486_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1494_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1502_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1510_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1518_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1526_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1534_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1542_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_154_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1550_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1558_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1566_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1574_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1582_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1590_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1598_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1606_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1614_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1622_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1630_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1638_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1646_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_164_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1654_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1662_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1670_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1678_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1686_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1694_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1702_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1710_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1718_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1726_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1734_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1742_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_174_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1750_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1758_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1766_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1774_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1782_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1790_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1798_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1806_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1814_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1822_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1830_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1838_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1846_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_184_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1854_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1862_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1870_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1878_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1886_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1894_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1902_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1910_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1918_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1926_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1934_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1942_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_194_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1950_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1958_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1966_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1974_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1982_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1990_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1998_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2006_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2014_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2022_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2030_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2038_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2046_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_204_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2054_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2062_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2070_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2078_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2086_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2094_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2102_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2110_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2118_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2126_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2134_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2142_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_214_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2150_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2158_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2166_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2174_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2182_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2190_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2198_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2206_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2214_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2222_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2230_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2238_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2246_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_224_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2254_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2262_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2270_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2278_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2286_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2294_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2302_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_234_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_244_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_24_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_254_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_264_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_274_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_284_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_294_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_304_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_314_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_324_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_334_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_344_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_34_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_354_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_364_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_374_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_384_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_394_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_404_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_414_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_424_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_434_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_444_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_44_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_454_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_464_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_474_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_484_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_494_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_504_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_514_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_524_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_534_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_544_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_54_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_554_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_564_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_574_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_584_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_594_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_604_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_614_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_624_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_634_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_644_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_64_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_654_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_664_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_674_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_684_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_694_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_704_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_714_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_724_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_734_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_744_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_74_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_754_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_764_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_774_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_784_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_794_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_804_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_814_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_824_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_834_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_844_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_84_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_854_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_864_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_874_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_884_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_894_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_904_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_914_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_924_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_934_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_944_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_94_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_954_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_964_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_974_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_984_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_994_wire : std_logic_vector(0 downto 0);
    signal IMA0_20 : std_logic_vector(7 downto 0);
    signal IMA100_1020 : std_logic_vector(7 downto 0);
    signal IMA101_1030 : std_logic_vector(7 downto 0);
    signal IMA102_1040 : std_logic_vector(7 downto 0);
    signal IMA103_1050 : std_logic_vector(7 downto 0);
    signal IMA104_1060 : std_logic_vector(7 downto 0);
    signal IMA105_1070 : std_logic_vector(7 downto 0);
    signal IMA106_1080 : std_logic_vector(7 downto 0);
    signal IMA107_1090 : std_logic_vector(7 downto 0);
    signal IMA108_1100 : std_logic_vector(7 downto 0);
    signal IMA109_1110 : std_logic_vector(7 downto 0);
    signal IMA10_120 : std_logic_vector(7 downto 0);
    signal IMA110_1120 : std_logic_vector(7 downto 0);
    signal IMA111_1130 : std_logic_vector(7 downto 0);
    signal IMA112_1140 : std_logic_vector(7 downto 0);
    signal IMA113_1150 : std_logic_vector(7 downto 0);
    signal IMA114_1160 : std_logic_vector(7 downto 0);
    signal IMA115_1170 : std_logic_vector(7 downto 0);
    signal IMA116_1180 : std_logic_vector(7 downto 0);
    signal IMA117_1190 : std_logic_vector(7 downto 0);
    signal IMA118_1200 : std_logic_vector(7 downto 0);
    signal IMA119_1210 : std_logic_vector(7 downto 0);
    signal IMA11_130 : std_logic_vector(7 downto 0);
    signal IMA120_1220 : std_logic_vector(7 downto 0);
    signal IMA121_1230 : std_logic_vector(7 downto 0);
    signal IMA122_1240 : std_logic_vector(7 downto 0);
    signal IMA123_1250 : std_logic_vector(7 downto 0);
    signal IMA124_1260 : std_logic_vector(7 downto 0);
    signal IMA125_1270 : std_logic_vector(7 downto 0);
    signal IMA126_1280 : std_logic_vector(7 downto 0);
    signal IMA127_1290 : std_logic_vector(7 downto 0);
    signal IMA12_140 : std_logic_vector(7 downto 0);
    signal IMA13_150 : std_logic_vector(7 downto 0);
    signal IMA14_160 : std_logic_vector(7 downto 0);
    signal IMA15_170 : std_logic_vector(7 downto 0);
    signal IMA16_180 : std_logic_vector(7 downto 0);
    signal IMA17_190 : std_logic_vector(7 downto 0);
    signal IMA18_200 : std_logic_vector(7 downto 0);
    signal IMA19_210 : std_logic_vector(7 downto 0);
    signal IMA1_30 : std_logic_vector(7 downto 0);
    signal IMA20_220 : std_logic_vector(7 downto 0);
    signal IMA21_230 : std_logic_vector(7 downto 0);
    signal IMA22_240 : std_logic_vector(7 downto 0);
    signal IMA23_250 : std_logic_vector(7 downto 0);
    signal IMA24_260 : std_logic_vector(7 downto 0);
    signal IMA25_270 : std_logic_vector(7 downto 0);
    signal IMA26_280 : std_logic_vector(7 downto 0);
    signal IMA27_290 : std_logic_vector(7 downto 0);
    signal IMA28_300 : std_logic_vector(7 downto 0);
    signal IMA29_310 : std_logic_vector(7 downto 0);
    signal IMA2_40 : std_logic_vector(7 downto 0);
    signal IMA30_320 : std_logic_vector(7 downto 0);
    signal IMA31_330 : std_logic_vector(7 downto 0);
    signal IMA32_340 : std_logic_vector(7 downto 0);
    signal IMA33_350 : std_logic_vector(7 downto 0);
    signal IMA34_360 : std_logic_vector(7 downto 0);
    signal IMA35_370 : std_logic_vector(7 downto 0);
    signal IMA36_380 : std_logic_vector(7 downto 0);
    signal IMA37_390 : std_logic_vector(7 downto 0);
    signal IMA38_400 : std_logic_vector(7 downto 0);
    signal IMA39_410 : std_logic_vector(7 downto 0);
    signal IMA3_50 : std_logic_vector(7 downto 0);
    signal IMA40_420 : std_logic_vector(7 downto 0);
    signal IMA41_430 : std_logic_vector(7 downto 0);
    signal IMA42_440 : std_logic_vector(7 downto 0);
    signal IMA43_450 : std_logic_vector(7 downto 0);
    signal IMA44_460 : std_logic_vector(7 downto 0);
    signal IMA45_470 : std_logic_vector(7 downto 0);
    signal IMA46_480 : std_logic_vector(7 downto 0);
    signal IMA47_490 : std_logic_vector(7 downto 0);
    signal IMA48_500 : std_logic_vector(7 downto 0);
    signal IMA49_510 : std_logic_vector(7 downto 0);
    signal IMA4_60 : std_logic_vector(7 downto 0);
    signal IMA50_520 : std_logic_vector(7 downto 0);
    signal IMA51_530 : std_logic_vector(7 downto 0);
    signal IMA52_540 : std_logic_vector(7 downto 0);
    signal IMA53_550 : std_logic_vector(7 downto 0);
    signal IMA54_560 : std_logic_vector(7 downto 0);
    signal IMA55_570 : std_logic_vector(7 downto 0);
    signal IMA56_580 : std_logic_vector(7 downto 0);
    signal IMA57_590 : std_logic_vector(7 downto 0);
    signal IMA58_600 : std_logic_vector(7 downto 0);
    signal IMA59_610 : std_logic_vector(7 downto 0);
    signal IMA5_70 : std_logic_vector(7 downto 0);
    signal IMA60_620 : std_logic_vector(7 downto 0);
    signal IMA61_630 : std_logic_vector(7 downto 0);
    signal IMA62_640 : std_logic_vector(7 downto 0);
    signal IMA63_650 : std_logic_vector(7 downto 0);
    signal IMA64_660 : std_logic_vector(7 downto 0);
    signal IMA65_670 : std_logic_vector(7 downto 0);
    signal IMA66_680 : std_logic_vector(7 downto 0);
    signal IMA67_690 : std_logic_vector(7 downto 0);
    signal IMA68_700 : std_logic_vector(7 downto 0);
    signal IMA69_710 : std_logic_vector(7 downto 0);
    signal IMA6_80 : std_logic_vector(7 downto 0);
    signal IMA70_720 : std_logic_vector(7 downto 0);
    signal IMA71_730 : std_logic_vector(7 downto 0);
    signal IMA72_740 : std_logic_vector(7 downto 0);
    signal IMA73_750 : std_logic_vector(7 downto 0);
    signal IMA74_760 : std_logic_vector(7 downto 0);
    signal IMA75_770 : std_logic_vector(7 downto 0);
    signal IMA76_780 : std_logic_vector(7 downto 0);
    signal IMA77_790 : std_logic_vector(7 downto 0);
    signal IMA78_800 : std_logic_vector(7 downto 0);
    signal IMA79_810 : std_logic_vector(7 downto 0);
    signal IMA7_90 : std_logic_vector(7 downto 0);
    signal IMA80_820 : std_logic_vector(7 downto 0);
    signal IMA81_830 : std_logic_vector(7 downto 0);
    signal IMA82_840 : std_logic_vector(7 downto 0);
    signal IMA83_850 : std_logic_vector(7 downto 0);
    signal IMA84_860 : std_logic_vector(7 downto 0);
    signal IMA85_870 : std_logic_vector(7 downto 0);
    signal IMA86_880 : std_logic_vector(7 downto 0);
    signal IMA87_890 : std_logic_vector(7 downto 0);
    signal IMA88_900 : std_logic_vector(7 downto 0);
    signal IMA89_910 : std_logic_vector(7 downto 0);
    signal IMA8_100 : std_logic_vector(7 downto 0);
    signal IMA90_920 : std_logic_vector(7 downto 0);
    signal IMA91_930 : std_logic_vector(7 downto 0);
    signal IMA92_940 : std_logic_vector(7 downto 0);
    signal IMA93_950 : std_logic_vector(7 downto 0);
    signal IMA94_960 : std_logic_vector(7 downto 0);
    signal IMA95_970 : std_logic_vector(7 downto 0);
    signal IMA96_980 : std_logic_vector(7 downto 0);
    signal IMA97_990 : std_logic_vector(7 downto 0);
    signal IMA98_1000 : std_logic_vector(7 downto 0);
    signal IMA99_1010 : std_logic_vector(7 downto 0);
    signal IMA9_110 : std_logic_vector(7 downto 0);
    signal IMB0_1298 : std_logic_vector(7 downto 0);
    signal IMB10_1378 : std_logic_vector(7 downto 0);
    signal IMB11_1386 : std_logic_vector(7 downto 0);
    signal IMB12_1394 : std_logic_vector(7 downto 0);
    signal IMB13_1402 : std_logic_vector(7 downto 0);
    signal IMB14_1410 : std_logic_vector(7 downto 0);
    signal IMB15_1418 : std_logic_vector(7 downto 0);
    signal IMB16_1426 : std_logic_vector(7 downto 0);
    signal IMB17_1434 : std_logic_vector(7 downto 0);
    signal IMB18_1442 : std_logic_vector(7 downto 0);
    signal IMB19_1450 : std_logic_vector(7 downto 0);
    signal IMB1_1306 : std_logic_vector(7 downto 0);
    signal IMB20_1458 : std_logic_vector(7 downto 0);
    signal IMB21_1466 : std_logic_vector(7 downto 0);
    signal IMB22_1474 : std_logic_vector(7 downto 0);
    signal IMB23_1482 : std_logic_vector(7 downto 0);
    signal IMB24_1490 : std_logic_vector(7 downto 0);
    signal IMB25_1498 : std_logic_vector(7 downto 0);
    signal IMB26_1506 : std_logic_vector(7 downto 0);
    signal IMB27_1514 : std_logic_vector(7 downto 0);
    signal IMB28_1522 : std_logic_vector(7 downto 0);
    signal IMB29_1530 : std_logic_vector(7 downto 0);
    signal IMB2_1314 : std_logic_vector(7 downto 0);
    signal IMB30_1538 : std_logic_vector(7 downto 0);
    signal IMB31_1546 : std_logic_vector(7 downto 0);
    signal IMB32_1554 : std_logic_vector(7 downto 0);
    signal IMB33_1562 : std_logic_vector(7 downto 0);
    signal IMB34_1570 : std_logic_vector(7 downto 0);
    signal IMB35_1578 : std_logic_vector(7 downto 0);
    signal IMB36_1586 : std_logic_vector(7 downto 0);
    signal IMB37_1594 : std_logic_vector(7 downto 0);
    signal IMB38_1602 : std_logic_vector(7 downto 0);
    signal IMB39_1610 : std_logic_vector(7 downto 0);
    signal IMB3_1322 : std_logic_vector(7 downto 0);
    signal IMB40_1618 : std_logic_vector(7 downto 0);
    signal IMB41_1626 : std_logic_vector(7 downto 0);
    signal IMB42_1634 : std_logic_vector(7 downto 0);
    signal IMB43_1642 : std_logic_vector(7 downto 0);
    signal IMB44_1650 : std_logic_vector(7 downto 0);
    signal IMB45_1658 : std_logic_vector(7 downto 0);
    signal IMB46_1666 : std_logic_vector(7 downto 0);
    signal IMB47_1674 : std_logic_vector(7 downto 0);
    signal IMB48_1682 : std_logic_vector(7 downto 0);
    signal IMB49_1690 : std_logic_vector(7 downto 0);
    signal IMB4_1330 : std_logic_vector(7 downto 0);
    signal IMB50_1698 : std_logic_vector(7 downto 0);
    signal IMB51_1706 : std_logic_vector(7 downto 0);
    signal IMB52_1714 : std_logic_vector(7 downto 0);
    signal IMB53_1722 : std_logic_vector(7 downto 0);
    signal IMB54_1730 : std_logic_vector(7 downto 0);
    signal IMB55_1738 : std_logic_vector(7 downto 0);
    signal IMB56_1746 : std_logic_vector(7 downto 0);
    signal IMB57_1754 : std_logic_vector(7 downto 0);
    signal IMB58_1762 : std_logic_vector(7 downto 0);
    signal IMB59_1770 : std_logic_vector(7 downto 0);
    signal IMB5_1338 : std_logic_vector(7 downto 0);
    signal IMB60_1778 : std_logic_vector(7 downto 0);
    signal IMB61_1786 : std_logic_vector(7 downto 0);
    signal IMB62_1794 : std_logic_vector(7 downto 0);
    signal IMB63_1802 : std_logic_vector(7 downto 0);
    signal IMB6_1346 : std_logic_vector(7 downto 0);
    signal IMB7_1354 : std_logic_vector(7 downto 0);
    signal IMB8_1362 : std_logic_vector(7 downto 0);
    signal IMB9_1370 : std_logic_vector(7 downto 0);
    signal IMC0_1810 : std_logic_vector(7 downto 0);
    signal IMC10_1890 : std_logic_vector(7 downto 0);
    signal IMC11_1898 : std_logic_vector(7 downto 0);
    signal IMC12_1906 : std_logic_vector(7 downto 0);
    signal IMC13_1914 : std_logic_vector(7 downto 0);
    signal IMC14_1922 : std_logic_vector(7 downto 0);
    signal IMC15_1930 : std_logic_vector(7 downto 0);
    signal IMC16_1938 : std_logic_vector(7 downto 0);
    signal IMC17_1946 : std_logic_vector(7 downto 0);
    signal IMC18_1954 : std_logic_vector(7 downto 0);
    signal IMC19_1962 : std_logic_vector(7 downto 0);
    signal IMC1_1818 : std_logic_vector(7 downto 0);
    signal IMC20_1970 : std_logic_vector(7 downto 0);
    signal IMC21_1978 : std_logic_vector(7 downto 0);
    signal IMC22_1986 : std_logic_vector(7 downto 0);
    signal IMC23_1994 : std_logic_vector(7 downto 0);
    signal IMC24_2002 : std_logic_vector(7 downto 0);
    signal IMC25_2010 : std_logic_vector(7 downto 0);
    signal IMC26_2018 : std_logic_vector(7 downto 0);
    signal IMC27_2026 : std_logic_vector(7 downto 0);
    signal IMC28_2034 : std_logic_vector(7 downto 0);
    signal IMC29_2042 : std_logic_vector(7 downto 0);
    signal IMC2_1826 : std_logic_vector(7 downto 0);
    signal IMC30_2050 : std_logic_vector(7 downto 0);
    signal IMC31_2058 : std_logic_vector(7 downto 0);
    signal IMC3_1834 : std_logic_vector(7 downto 0);
    signal IMC4_1842 : std_logic_vector(7 downto 0);
    signal IMC5_1850 : std_logic_vector(7 downto 0);
    signal IMC6_1858 : std_logic_vector(7 downto 0);
    signal IMC7_1866 : std_logic_vector(7 downto 0);
    signal IMC8_1874 : std_logic_vector(7 downto 0);
    signal IMC9_1882 : std_logic_vector(7 downto 0);
    signal IMD0_2066 : std_logic_vector(7 downto 0);
    signal IMD10_2146 : std_logic_vector(7 downto 0);
    signal IMD11_2154 : std_logic_vector(7 downto 0);
    signal IMD12_2162 : std_logic_vector(7 downto 0);
    signal IMD13_2170 : std_logic_vector(7 downto 0);
    signal IMD14_2178 : std_logic_vector(7 downto 0);
    signal IMD15_2186 : std_logic_vector(7 downto 0);
    signal IMD1_2074 : std_logic_vector(7 downto 0);
    signal IMD2_2082 : std_logic_vector(7 downto 0);
    signal IMD3_2090 : std_logic_vector(7 downto 0);
    signal IMD4_2098 : std_logic_vector(7 downto 0);
    signal IMD5_2106 : std_logic_vector(7 downto 0);
    signal IMD6_2114 : std_logic_vector(7 downto 0);
    signal IMD7_2122 : std_logic_vector(7 downto 0);
    signal IMD8_2130 : std_logic_vector(7 downto 0);
    signal IMD9_2138 : std_logic_vector(7 downto 0);
    signal IME0_2194 : std_logic_vector(7 downto 0);
    signal IME1_2202 : std_logic_vector(7 downto 0);
    signal IME2_2210 : std_logic_vector(7 downto 0);
    signal IME3_2218 : std_logic_vector(7 downto 0);
    signal IME4_2226 : std_logic_vector(7 downto 0);
    signal IME5_2234 : std_logic_vector(7 downto 0);
    signal IME6_2242 : std_logic_vector(7 downto 0);
    signal IME7_2250 : std_logic_vector(7 downto 0);
    signal IMF0_2258 : std_logic_vector(7 downto 0);
    signal IMF1_2266 : std_logic_vector(7 downto 0);
    signal IMF2_2274 : std_logic_vector(7 downto 0);
    signal IMF3_2282 : std_logic_vector(7 downto 0);
    signal IMG0_2290 : std_logic_vector(7 downto 0);
    signal IMG1_2298 : std_logic_vector(7 downto 0);
    signal konst_1003_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1013_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1023_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1033_wire_constant : std_logic_vector(7 downto 0);
    signal konst_103_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1043_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1053_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1063_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1073_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1083_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1093_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1103_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1113_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1123_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1133_wire_constant : std_logic_vector(7 downto 0);
    signal konst_113_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1143_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1153_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1163_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1173_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1183_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1193_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1203_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1213_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1223_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1233_wire_constant : std_logic_vector(7 downto 0);
    signal konst_123_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1243_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1253_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1263_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1273_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1283_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1293_wire_constant : std_logic_vector(7 downto 0);
    signal konst_12_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1301_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1309_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1317_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1325_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1333_wire_constant : std_logic_vector(7 downto 0);
    signal konst_133_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1341_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1349_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1357_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1365_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1373_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1381_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1389_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1397_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1405_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1413_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1421_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1429_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1437_wire_constant : std_logic_vector(7 downto 0);
    signal konst_143_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1445_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1453_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1461_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1469_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1477_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1485_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1493_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1501_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1509_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1517_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1525_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1533_wire_constant : std_logic_vector(7 downto 0);
    signal konst_153_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1541_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1549_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1557_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1565_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1573_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1581_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1589_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1597_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1605_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1613_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1621_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1629_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1637_wire_constant : std_logic_vector(7 downto 0);
    signal konst_163_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1645_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1653_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1661_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1669_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1677_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1685_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1693_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1701_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1709_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1717_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1725_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1733_wire_constant : std_logic_vector(7 downto 0);
    signal konst_173_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1741_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1749_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1757_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1765_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1773_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1781_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1789_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1797_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1805_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1813_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1821_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1829_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1837_wire_constant : std_logic_vector(7 downto 0);
    signal konst_183_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1845_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1853_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1861_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1869_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1877_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1885_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1893_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1901_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1909_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1917_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1925_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1933_wire_constant : std_logic_vector(7 downto 0);
    signal konst_193_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1941_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1949_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1957_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1965_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1973_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1981_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1989_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1997_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2005_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2013_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2021_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2029_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2037_wire_constant : std_logic_vector(7 downto 0);
    signal konst_203_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2045_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2053_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2061_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2069_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2077_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2085_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2093_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2101_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2109_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2117_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2125_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2133_wire_constant : std_logic_vector(7 downto 0);
    signal konst_213_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2141_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2149_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2157_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2165_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2173_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2181_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2189_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2197_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2205_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2213_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2221_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2229_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2237_wire_constant : std_logic_vector(7 downto 0);
    signal konst_223_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2245_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2253_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2261_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2269_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2277_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2285_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2293_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2301_wire_constant : std_logic_vector(7 downto 0);
    signal konst_233_wire_constant : std_logic_vector(7 downto 0);
    signal konst_23_wire_constant : std_logic_vector(7 downto 0);
    signal konst_243_wire_constant : std_logic_vector(7 downto 0);
    signal konst_253_wire_constant : std_logic_vector(7 downto 0);
    signal konst_263_wire_constant : std_logic_vector(7 downto 0);
    signal konst_273_wire_constant : std_logic_vector(7 downto 0);
    signal konst_283_wire_constant : std_logic_vector(7 downto 0);
    signal konst_293_wire_constant : std_logic_vector(7 downto 0);
    signal konst_303_wire_constant : std_logic_vector(7 downto 0);
    signal konst_313_wire_constant : std_logic_vector(7 downto 0);
    signal konst_323_wire_constant : std_logic_vector(7 downto 0);
    signal konst_333_wire_constant : std_logic_vector(7 downto 0);
    signal konst_33_wire_constant : std_logic_vector(7 downto 0);
    signal konst_343_wire_constant : std_logic_vector(7 downto 0);
    signal konst_353_wire_constant : std_logic_vector(7 downto 0);
    signal konst_363_wire_constant : std_logic_vector(7 downto 0);
    signal konst_373_wire_constant : std_logic_vector(7 downto 0);
    signal konst_383_wire_constant : std_logic_vector(7 downto 0);
    signal konst_393_wire_constant : std_logic_vector(7 downto 0);
    signal konst_403_wire_constant : std_logic_vector(7 downto 0);
    signal konst_413_wire_constant : std_logic_vector(7 downto 0);
    signal konst_423_wire_constant : std_logic_vector(7 downto 0);
    signal konst_433_wire_constant : std_logic_vector(7 downto 0);
    signal konst_43_wire_constant : std_logic_vector(7 downto 0);
    signal konst_443_wire_constant : std_logic_vector(7 downto 0);
    signal konst_453_wire_constant : std_logic_vector(7 downto 0);
    signal konst_463_wire_constant : std_logic_vector(7 downto 0);
    signal konst_473_wire_constant : std_logic_vector(7 downto 0);
    signal konst_483_wire_constant : std_logic_vector(7 downto 0);
    signal konst_493_wire_constant : std_logic_vector(7 downto 0);
    signal konst_503_wire_constant : std_logic_vector(7 downto 0);
    signal konst_513_wire_constant : std_logic_vector(7 downto 0);
    signal konst_523_wire_constant : std_logic_vector(7 downto 0);
    signal konst_533_wire_constant : std_logic_vector(7 downto 0);
    signal konst_53_wire_constant : std_logic_vector(7 downto 0);
    signal konst_543_wire_constant : std_logic_vector(7 downto 0);
    signal konst_553_wire_constant : std_logic_vector(7 downto 0);
    signal konst_563_wire_constant : std_logic_vector(7 downto 0);
    signal konst_573_wire_constant : std_logic_vector(7 downto 0);
    signal konst_583_wire_constant : std_logic_vector(7 downto 0);
    signal konst_593_wire_constant : std_logic_vector(7 downto 0);
    signal konst_603_wire_constant : std_logic_vector(7 downto 0);
    signal konst_613_wire_constant : std_logic_vector(7 downto 0);
    signal konst_623_wire_constant : std_logic_vector(7 downto 0);
    signal konst_633_wire_constant : std_logic_vector(7 downto 0);
    signal konst_63_wire_constant : std_logic_vector(7 downto 0);
    signal konst_643_wire_constant : std_logic_vector(7 downto 0);
    signal konst_653_wire_constant : std_logic_vector(7 downto 0);
    signal konst_663_wire_constant : std_logic_vector(7 downto 0);
    signal konst_673_wire_constant : std_logic_vector(7 downto 0);
    signal konst_683_wire_constant : std_logic_vector(7 downto 0);
    signal konst_693_wire_constant : std_logic_vector(7 downto 0);
    signal konst_703_wire_constant : std_logic_vector(7 downto 0);
    signal konst_713_wire_constant : std_logic_vector(7 downto 0);
    signal konst_723_wire_constant : std_logic_vector(7 downto 0);
    signal konst_733_wire_constant : std_logic_vector(7 downto 0);
    signal konst_73_wire_constant : std_logic_vector(7 downto 0);
    signal konst_743_wire_constant : std_logic_vector(7 downto 0);
    signal konst_753_wire_constant : std_logic_vector(7 downto 0);
    signal konst_763_wire_constant : std_logic_vector(7 downto 0);
    signal konst_773_wire_constant : std_logic_vector(7 downto 0);
    signal konst_783_wire_constant : std_logic_vector(7 downto 0);
    signal konst_793_wire_constant : std_logic_vector(7 downto 0);
    signal konst_803_wire_constant : std_logic_vector(7 downto 0);
    signal konst_813_wire_constant : std_logic_vector(7 downto 0);
    signal konst_823_wire_constant : std_logic_vector(7 downto 0);
    signal konst_833_wire_constant : std_logic_vector(7 downto 0);
    signal konst_83_wire_constant : std_logic_vector(7 downto 0);
    signal konst_843_wire_constant : std_logic_vector(7 downto 0);
    signal konst_853_wire_constant : std_logic_vector(7 downto 0);
    signal konst_863_wire_constant : std_logic_vector(7 downto 0);
    signal konst_873_wire_constant : std_logic_vector(7 downto 0);
    signal konst_883_wire_constant : std_logic_vector(7 downto 0);
    signal konst_893_wire_constant : std_logic_vector(7 downto 0);
    signal konst_903_wire_constant : std_logic_vector(7 downto 0);
    signal konst_913_wire_constant : std_logic_vector(7 downto 0);
    signal konst_923_wire_constant : std_logic_vector(7 downto 0);
    signal konst_933_wire_constant : std_logic_vector(7 downto 0);
    signal konst_93_wire_constant : std_logic_vector(7 downto 0);
    signal konst_943_wire_constant : std_logic_vector(7 downto 0);
    signal konst_953_wire_constant : std_logic_vector(7 downto 0);
    signal konst_963_wire_constant : std_logic_vector(7 downto 0);
    signal konst_973_wire_constant : std_logic_vector(7 downto 0);
    signal konst_983_wire_constant : std_logic_vector(7 downto 0);
    signal konst_993_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1006_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1008_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1016_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1018_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1026_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1028_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1036_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1038_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1046_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1048_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1056_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1058_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1066_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1068_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_106_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1076_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1078_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1086_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1088_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_108_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1096_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1098_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1106_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1108_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1116_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1118_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1126_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1128_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1136_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1138_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1146_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1148_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1156_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1158_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1166_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1168_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_116_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1176_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1178_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1186_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1188_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_118_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1196_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1198_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1206_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1208_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1216_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1218_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1226_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1228_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1236_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1238_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1246_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1248_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1256_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1258_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1266_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1268_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_126_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1276_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1278_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1286_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1288_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_128_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_136_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_138_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_146_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_148_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_156_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_158_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_166_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_168_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_16_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_176_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_178_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_186_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_188_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_18_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_196_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_198_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_206_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_208_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_216_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_218_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_226_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_228_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_236_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_238_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_246_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_248_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_256_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_258_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_266_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_268_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_26_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_276_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_278_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_286_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_288_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_28_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_296_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_298_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_306_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_308_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_316_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_318_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_326_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_328_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_336_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_338_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_346_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_348_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_356_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_358_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_366_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_368_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_36_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_376_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_378_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_386_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_388_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_38_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_396_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_398_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_406_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_408_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_416_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_418_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_426_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_428_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_436_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_438_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_446_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_448_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_456_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_458_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_466_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_468_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_46_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_476_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_478_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_486_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_488_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_48_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_496_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_498_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_506_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_508_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_516_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_518_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_526_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_528_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_536_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_538_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_546_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_548_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_556_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_558_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_566_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_568_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_56_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_576_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_578_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_586_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_588_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_58_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_596_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_598_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_606_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_608_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_616_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_618_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_626_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_628_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_636_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_638_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_646_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_648_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_656_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_658_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_666_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_668_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_66_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_676_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_678_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_686_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_688_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_68_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_696_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_698_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_706_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_708_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_716_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_718_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_726_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_728_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_736_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_738_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_746_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_748_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_756_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_758_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_766_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_768_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_76_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_776_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_778_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_786_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_788_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_78_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_796_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_798_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_806_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_808_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_816_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_818_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_826_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_828_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_836_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_838_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_846_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_848_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_856_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_858_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_866_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_868_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_86_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_876_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_878_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_886_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_888_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_88_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_896_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_898_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_906_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_908_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_916_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_918_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_926_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_928_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_936_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_938_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_946_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_948_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_956_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_958_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_966_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_968_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_96_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_976_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_978_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_986_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_988_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_98_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_996_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_998_wire_constant : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    konst_1003_wire_constant <= "00000000";
    konst_1013_wire_constant <= "00000000";
    konst_1023_wire_constant <= "00000000";
    konst_1033_wire_constant <= "00000000";
    konst_103_wire_constant <= "00000000";
    konst_1043_wire_constant <= "00000000";
    konst_1053_wire_constant <= "00000000";
    konst_1063_wire_constant <= "00000000";
    konst_1073_wire_constant <= "00000000";
    konst_1083_wire_constant <= "00000000";
    konst_1093_wire_constant <= "00000000";
    konst_1103_wire_constant <= "00000000";
    konst_1113_wire_constant <= "00000000";
    konst_1123_wire_constant <= "00000000";
    konst_1133_wire_constant <= "00000000";
    konst_113_wire_constant <= "00000000";
    konst_1143_wire_constant <= "00000000";
    konst_1153_wire_constant <= "00000000";
    konst_1163_wire_constant <= "00000000";
    konst_1173_wire_constant <= "00000000";
    konst_1183_wire_constant <= "00000000";
    konst_1193_wire_constant <= "00000000";
    konst_1203_wire_constant <= "00000000";
    konst_1213_wire_constant <= "00000000";
    konst_1223_wire_constant <= "00000000";
    konst_1233_wire_constant <= "00000000";
    konst_123_wire_constant <= "00000000";
    konst_1243_wire_constant <= "00000000";
    konst_1253_wire_constant <= "00000000";
    konst_1263_wire_constant <= "00000000";
    konst_1273_wire_constant <= "00000000";
    konst_1283_wire_constant <= "00000000";
    konst_1293_wire_constant <= "00000001";
    konst_12_wire_constant <= "00000000";
    konst_1301_wire_constant <= "00000001";
    konst_1309_wire_constant <= "00000001";
    konst_1317_wire_constant <= "00000001";
    konst_1325_wire_constant <= "00000001";
    konst_1333_wire_constant <= "00000001";
    konst_133_wire_constant <= "00000000";
    konst_1341_wire_constant <= "00000001";
    konst_1349_wire_constant <= "00000001";
    konst_1357_wire_constant <= "00000001";
    konst_1365_wire_constant <= "00000001";
    konst_1373_wire_constant <= "00000001";
    konst_1381_wire_constant <= "00000001";
    konst_1389_wire_constant <= "00000001";
    konst_1397_wire_constant <= "00000001";
    konst_1405_wire_constant <= "00000001";
    konst_1413_wire_constant <= "00000001";
    konst_1421_wire_constant <= "00000001";
    konst_1429_wire_constant <= "00000001";
    konst_1437_wire_constant <= "00000001";
    konst_143_wire_constant <= "00000000";
    konst_1445_wire_constant <= "00000001";
    konst_1453_wire_constant <= "00000001";
    konst_1461_wire_constant <= "00000001";
    konst_1469_wire_constant <= "00000001";
    konst_1477_wire_constant <= "00000001";
    konst_1485_wire_constant <= "00000001";
    konst_1493_wire_constant <= "00000001";
    konst_1501_wire_constant <= "00000001";
    konst_1509_wire_constant <= "00000001";
    konst_1517_wire_constant <= "00000001";
    konst_1525_wire_constant <= "00000001";
    konst_1533_wire_constant <= "00000001";
    konst_153_wire_constant <= "00000000";
    konst_1541_wire_constant <= "00000001";
    konst_1549_wire_constant <= "00000001";
    konst_1557_wire_constant <= "00000001";
    konst_1565_wire_constant <= "00000001";
    konst_1573_wire_constant <= "00000001";
    konst_1581_wire_constant <= "00000001";
    konst_1589_wire_constant <= "00000001";
    konst_1597_wire_constant <= "00000001";
    konst_1605_wire_constant <= "00000001";
    konst_1613_wire_constant <= "00000001";
    konst_1621_wire_constant <= "00000001";
    konst_1629_wire_constant <= "00000001";
    konst_1637_wire_constant <= "00000001";
    konst_163_wire_constant <= "00000000";
    konst_1645_wire_constant <= "00000001";
    konst_1653_wire_constant <= "00000001";
    konst_1661_wire_constant <= "00000001";
    konst_1669_wire_constant <= "00000001";
    konst_1677_wire_constant <= "00000001";
    konst_1685_wire_constant <= "00000001";
    konst_1693_wire_constant <= "00000001";
    konst_1701_wire_constant <= "00000001";
    konst_1709_wire_constant <= "00000001";
    konst_1717_wire_constant <= "00000001";
    konst_1725_wire_constant <= "00000001";
    konst_1733_wire_constant <= "00000001";
    konst_173_wire_constant <= "00000000";
    konst_1741_wire_constant <= "00000001";
    konst_1749_wire_constant <= "00000001";
    konst_1757_wire_constant <= "00000001";
    konst_1765_wire_constant <= "00000001";
    konst_1773_wire_constant <= "00000001";
    konst_1781_wire_constant <= "00000001";
    konst_1789_wire_constant <= "00000001";
    konst_1797_wire_constant <= "00000001";
    konst_1805_wire_constant <= "00000010";
    konst_1813_wire_constant <= "00000010";
    konst_1821_wire_constant <= "00000010";
    konst_1829_wire_constant <= "00000010";
    konst_1837_wire_constant <= "00000010";
    konst_183_wire_constant <= "00000000";
    konst_1845_wire_constant <= "00000010";
    konst_1853_wire_constant <= "00000010";
    konst_1861_wire_constant <= "00000010";
    konst_1869_wire_constant <= "00000010";
    konst_1877_wire_constant <= "00000010";
    konst_1885_wire_constant <= "00000010";
    konst_1893_wire_constant <= "00000010";
    konst_1901_wire_constant <= "00000010";
    konst_1909_wire_constant <= "00000010";
    konst_1917_wire_constant <= "00000010";
    konst_1925_wire_constant <= "00000010";
    konst_1933_wire_constant <= "00000010";
    konst_193_wire_constant <= "00000000";
    konst_1941_wire_constant <= "00000010";
    konst_1949_wire_constant <= "00000010";
    konst_1957_wire_constant <= "00000010";
    konst_1965_wire_constant <= "00000010";
    konst_1973_wire_constant <= "00000010";
    konst_1981_wire_constant <= "00000010";
    konst_1989_wire_constant <= "00000010";
    konst_1997_wire_constant <= "00000010";
    konst_2005_wire_constant <= "00000010";
    konst_2013_wire_constant <= "00000010";
    konst_2021_wire_constant <= "00000010";
    konst_2029_wire_constant <= "00000010";
    konst_2037_wire_constant <= "00000010";
    konst_203_wire_constant <= "00000000";
    konst_2045_wire_constant <= "00000010";
    konst_2053_wire_constant <= "00000010";
    konst_2061_wire_constant <= "00000011";
    konst_2069_wire_constant <= "00000011";
    konst_2077_wire_constant <= "00000011";
    konst_2085_wire_constant <= "00000011";
    konst_2093_wire_constant <= "00000011";
    konst_2101_wire_constant <= "00000011";
    konst_2109_wire_constant <= "00000011";
    konst_2117_wire_constant <= "00000011";
    konst_2125_wire_constant <= "00000011";
    konst_2133_wire_constant <= "00000011";
    konst_213_wire_constant <= "00000000";
    konst_2141_wire_constant <= "00000011";
    konst_2149_wire_constant <= "00000011";
    konst_2157_wire_constant <= "00000011";
    konst_2165_wire_constant <= "00000011";
    konst_2173_wire_constant <= "00000011";
    konst_2181_wire_constant <= "00000011";
    konst_2189_wire_constant <= "00000100";
    konst_2197_wire_constant <= "00000100";
    konst_2205_wire_constant <= "00000100";
    konst_2213_wire_constant <= "00000100";
    konst_2221_wire_constant <= "00000100";
    konst_2229_wire_constant <= "00000100";
    konst_2237_wire_constant <= "00000100";
    konst_223_wire_constant <= "00000000";
    konst_2245_wire_constant <= "00000100";
    konst_2253_wire_constant <= "00000101";
    konst_2261_wire_constant <= "00000101";
    konst_2269_wire_constant <= "00000101";
    konst_2277_wire_constant <= "00000101";
    konst_2285_wire_constant <= "00000110";
    konst_2293_wire_constant <= "00000110";
    konst_2301_wire_constant <= "00000111";
    konst_233_wire_constant <= "00000000";
    konst_23_wire_constant <= "00000000";
    konst_243_wire_constant <= "00000000";
    konst_253_wire_constant <= "00000000";
    konst_263_wire_constant <= "00000000";
    konst_273_wire_constant <= "00000000";
    konst_283_wire_constant <= "00000000";
    konst_293_wire_constant <= "00000000";
    konst_303_wire_constant <= "00000000";
    konst_313_wire_constant <= "00000000";
    konst_323_wire_constant <= "00000000";
    konst_333_wire_constant <= "00000000";
    konst_33_wire_constant <= "00000000";
    konst_343_wire_constant <= "00000000";
    konst_353_wire_constant <= "00000000";
    konst_363_wire_constant <= "00000000";
    konst_373_wire_constant <= "00000000";
    konst_383_wire_constant <= "00000000";
    konst_393_wire_constant <= "00000000";
    konst_403_wire_constant <= "00000000";
    konst_413_wire_constant <= "00000000";
    konst_423_wire_constant <= "00000000";
    konst_433_wire_constant <= "00000000";
    konst_43_wire_constant <= "00000000";
    konst_443_wire_constant <= "00000000";
    konst_453_wire_constant <= "00000000";
    konst_463_wire_constant <= "00000000";
    konst_473_wire_constant <= "00000000";
    konst_483_wire_constant <= "00000000";
    konst_493_wire_constant <= "00000000";
    konst_503_wire_constant <= "00000000";
    konst_513_wire_constant <= "00000000";
    konst_523_wire_constant <= "00000000";
    konst_533_wire_constant <= "00000000";
    konst_53_wire_constant <= "00000000";
    konst_543_wire_constant <= "00000000";
    konst_553_wire_constant <= "00000000";
    konst_563_wire_constant <= "00000000";
    konst_573_wire_constant <= "00000000";
    konst_583_wire_constant <= "00000000";
    konst_593_wire_constant <= "00000000";
    konst_603_wire_constant <= "00000000";
    konst_613_wire_constant <= "00000000";
    konst_623_wire_constant <= "00000000";
    konst_633_wire_constant <= "00000000";
    konst_63_wire_constant <= "00000000";
    konst_643_wire_constant <= "00000000";
    konst_653_wire_constant <= "00000000";
    konst_663_wire_constant <= "00000000";
    konst_673_wire_constant <= "00000000";
    konst_683_wire_constant <= "00000000";
    konst_693_wire_constant <= "00000000";
    konst_703_wire_constant <= "00000000";
    konst_713_wire_constant <= "00000000";
    konst_723_wire_constant <= "00000000";
    konst_733_wire_constant <= "00000000";
    konst_73_wire_constant <= "00000000";
    konst_743_wire_constant <= "00000000";
    konst_753_wire_constant <= "00000000";
    konst_763_wire_constant <= "00000000";
    konst_773_wire_constant <= "00000000";
    konst_783_wire_constant <= "00000000";
    konst_793_wire_constant <= "00000000";
    konst_803_wire_constant <= "00000000";
    konst_813_wire_constant <= "00000000";
    konst_823_wire_constant <= "00000000";
    konst_833_wire_constant <= "00000000";
    konst_83_wire_constant <= "00000000";
    konst_843_wire_constant <= "00000000";
    konst_853_wire_constant <= "00000000";
    konst_863_wire_constant <= "00000000";
    konst_873_wire_constant <= "00000000";
    konst_883_wire_constant <= "00000000";
    konst_893_wire_constant <= "00000000";
    konst_903_wire_constant <= "00000000";
    konst_913_wire_constant <= "00000000";
    konst_923_wire_constant <= "00000000";
    konst_933_wire_constant <= "00000000";
    konst_93_wire_constant <= "00000000";
    konst_943_wire_constant <= "00000000";
    konst_953_wire_constant <= "00000000";
    konst_963_wire_constant <= "00000000";
    konst_973_wire_constant <= "00000000";
    konst_983_wire_constant <= "00000000";
    konst_993_wire_constant <= "00000000";
    type_cast_1006_wire_constant <= "00110001";
    type_cast_1008_wire_constant <= "11000111";
    type_cast_1016_wire_constant <= "00010010";
    type_cast_1018_wire_constant <= "10110001";
    type_cast_1026_wire_constant <= "01011001";
    type_cast_1028_wire_constant <= "00010000";
    type_cast_1036_wire_constant <= "10000000";
    type_cast_1038_wire_constant <= "00100111";
    type_cast_1046_wire_constant <= "01011111";
    type_cast_1048_wire_constant <= "11101100";
    type_cast_1056_wire_constant <= "01010001";
    type_cast_1058_wire_constant <= "01100000";
    type_cast_1066_wire_constant <= "10101001";
    type_cast_1068_wire_constant <= "01111111";
    type_cast_106_wire_constant <= "10000010";
    type_cast_1076_wire_constant <= "10110101";
    type_cast_1078_wire_constant <= "00011001";
    type_cast_1086_wire_constant <= "00001101";
    type_cast_1088_wire_constant <= "01001010";
    type_cast_108_wire_constant <= "00111001";
    type_cast_1096_wire_constant <= "11100101";
    type_cast_1098_wire_constant <= "00101101";
    type_cast_1106_wire_constant <= "10011111";
    type_cast_1108_wire_constant <= "01111010";
    type_cast_1116_wire_constant <= "11001001";
    type_cast_1118_wire_constant <= "10010011";
    type_cast_1126_wire_constant <= "11101111";
    type_cast_1128_wire_constant <= "10011100";
    type_cast_1136_wire_constant <= "11100000";
    type_cast_1138_wire_constant <= "10100000";
    type_cast_1146_wire_constant <= "01001101";
    type_cast_1148_wire_constant <= "00111011";
    type_cast_1156_wire_constant <= "00101010";
    type_cast_1158_wire_constant <= "10101110";
    type_cast_1166_wire_constant <= "10110000";
    type_cast_1168_wire_constant <= "11110101";
    type_cast_116_wire_constant <= "00101111";
    type_cast_1176_wire_constant <= "11101011";
    type_cast_1178_wire_constant <= "11001000";
    type_cast_1186_wire_constant <= "00111100";
    type_cast_1188_wire_constant <= "10111011";
    type_cast_118_wire_constant <= "10011011";
    type_cast_1196_wire_constant <= "01010011";
    type_cast_1198_wire_constant <= "10000011";
    type_cast_1206_wire_constant <= "01100001";
    type_cast_1208_wire_constant <= "10011001";
    type_cast_1216_wire_constant <= "00101011";
    type_cast_1218_wire_constant <= "00010111";
    type_cast_1226_wire_constant <= "01111110";
    type_cast_1228_wire_constant <= "00000100";
    type_cast_1236_wire_constant <= "01110111";
    type_cast_1238_wire_constant <= "10111010";
    type_cast_1246_wire_constant <= "00100110";
    type_cast_1248_wire_constant <= "11010110";
    type_cast_1256_wire_constant <= "01101001";
    type_cast_1258_wire_constant <= "11100001";
    type_cast_1266_wire_constant <= "01100011";
    type_cast_1268_wire_constant <= "00010100";
    type_cast_126_wire_constant <= "10000111";
    type_cast_1276_wire_constant <= "00100001";
    type_cast_1278_wire_constant <= "01010101";
    type_cast_1286_wire_constant <= "01111101";
    type_cast_1288_wire_constant <= "00001100";
    type_cast_128_wire_constant <= "11111111";
    type_cast_136_wire_constant <= "10001110";
    type_cast_138_wire_constant <= "00110100";
    type_cast_146_wire_constant <= "01000100";
    type_cast_148_wire_constant <= "01000011";
    type_cast_156_wire_constant <= "11011110";
    type_cast_158_wire_constant <= "11000100";
    type_cast_166_wire_constant <= "11001011";
    type_cast_168_wire_constant <= "11101001";
    type_cast_16_wire_constant <= "00001001";
    type_cast_176_wire_constant <= "01111011";
    type_cast_178_wire_constant <= "01010100";
    type_cast_186_wire_constant <= "00110010";
    type_cast_188_wire_constant <= "10010100";
    type_cast_18_wire_constant <= "01010010";
    type_cast_196_wire_constant <= "11000010";
    type_cast_198_wire_constant <= "10100110";
    type_cast_206_wire_constant <= "00111101";
    type_cast_208_wire_constant <= "00100011";
    type_cast_216_wire_constant <= "01001100";
    type_cast_218_wire_constant <= "11101110";
    type_cast_226_wire_constant <= "00001011";
    type_cast_228_wire_constant <= "10010101";
    type_cast_236_wire_constant <= "11111010";
    type_cast_238_wire_constant <= "01000010";
    type_cast_246_wire_constant <= "01001110";
    type_cast_248_wire_constant <= "11000011";
    type_cast_256_wire_constant <= "00101110";
    type_cast_258_wire_constant <= "00001000";
    type_cast_266_wire_constant <= "01100110";
    type_cast_268_wire_constant <= "10100001";
    type_cast_26_wire_constant <= "11010101";
    type_cast_276_wire_constant <= "11011001";
    type_cast_278_wire_constant <= "00101000";
    type_cast_286_wire_constant <= "10110010";
    type_cast_288_wire_constant <= "00100100";
    type_cast_28_wire_constant <= "01101010";
    type_cast_296_wire_constant <= "01011011";
    type_cast_298_wire_constant <= "01110110";
    type_cast_306_wire_constant <= "01001001";
    type_cast_308_wire_constant <= "10100010";
    type_cast_316_wire_constant <= "10001011";
    type_cast_318_wire_constant <= "01101101";
    type_cast_326_wire_constant <= "00100101";
    type_cast_328_wire_constant <= "11010001";
    type_cast_336_wire_constant <= "11111000";
    type_cast_338_wire_constant <= "01110010";
    type_cast_346_wire_constant <= "01100100";
    type_cast_348_wire_constant <= "11110110";
    type_cast_356_wire_constant <= "01101000";
    type_cast_358_wire_constant <= "10000110";
    type_cast_366_wire_constant <= "00010110";
    type_cast_368_wire_constant <= "10011000";
    type_cast_36_wire_constant <= "00110110";
    type_cast_376_wire_constant <= "10100100";
    type_cast_378_wire_constant <= "11010100";
    type_cast_386_wire_constant <= "11001100";
    type_cast_388_wire_constant <= "01011100";
    type_cast_38_wire_constant <= "00110000";
    type_cast_396_wire_constant <= "01100101";
    type_cast_398_wire_constant <= "01011101";
    type_cast_406_wire_constant <= "10010010";
    type_cast_408_wire_constant <= "10110110";
    type_cast_416_wire_constant <= "01110000";
    type_cast_418_wire_constant <= "01101100";
    type_cast_426_wire_constant <= "01010000";
    type_cast_428_wire_constant <= "01001000";
    type_cast_436_wire_constant <= "11101101";
    type_cast_438_wire_constant <= "11111101";
    type_cast_446_wire_constant <= "11011010";
    type_cast_448_wire_constant <= "10111001";
    type_cast_456_wire_constant <= "00010101";
    type_cast_458_wire_constant <= "01011110";
    type_cast_466_wire_constant <= "01010111";
    type_cast_468_wire_constant <= "01000110";
    type_cast_46_wire_constant <= "00111000";
    type_cast_476_wire_constant <= "10001101";
    type_cast_478_wire_constant <= "10100111";
    type_cast_486_wire_constant <= "10000100";
    type_cast_488_wire_constant <= "10011101";
    type_cast_48_wire_constant <= "10100101";
    type_cast_496_wire_constant <= "11011000";
    type_cast_498_wire_constant <= "10010000";
    type_cast_506_wire_constant <= "00000000";
    type_cast_508_wire_constant <= "10101011";
    type_cast_516_wire_constant <= "10111100";
    type_cast_518_wire_constant <= "10001100";
    type_cast_526_wire_constant <= "00001010";
    type_cast_528_wire_constant <= "11010011";
    type_cast_536_wire_constant <= "11100100";
    type_cast_538_wire_constant <= "11110111";
    type_cast_546_wire_constant <= "00000101";
    type_cast_548_wire_constant <= "01011000";
    type_cast_556_wire_constant <= "10110011";
    type_cast_558_wire_constant <= "10111000";
    type_cast_566_wire_constant <= "00000110";
    type_cast_568_wire_constant <= "01000101";
    type_cast_56_wire_constant <= "01000000";
    type_cast_576_wire_constant <= "00101100";
    type_cast_578_wire_constant <= "11010000";
    type_cast_586_wire_constant <= "10001111";
    type_cast_588_wire_constant <= "00011110";
    type_cast_58_wire_constant <= "10111111";
    type_cast_596_wire_constant <= "00111111";
    type_cast_598_wire_constant <= "11001010";
    type_cast_606_wire_constant <= "00000010";
    type_cast_608_wire_constant <= "00001111";
    type_cast_616_wire_constant <= "10101111";
    type_cast_618_wire_constant <= "11000001";
    type_cast_626_wire_constant <= "00000011";
    type_cast_628_wire_constant <= "10111101";
    type_cast_636_wire_constant <= "00010011";
    type_cast_638_wire_constant <= "00000001";
    type_cast_646_wire_constant <= "01101011";
    type_cast_648_wire_constant <= "10001010";
    type_cast_656_wire_constant <= "10010001";
    type_cast_658_wire_constant <= "00111010";
    type_cast_666_wire_constant <= "01000001";
    type_cast_668_wire_constant <= "00010001";
    type_cast_66_wire_constant <= "10011110";
    type_cast_676_wire_constant <= "01100111";
    type_cast_678_wire_constant <= "01001111";
    type_cast_686_wire_constant <= "11101010";
    type_cast_688_wire_constant <= "11011100";
    type_cast_68_wire_constant <= "10100011";
    type_cast_696_wire_constant <= "11110010";
    type_cast_698_wire_constant <= "10010111";
    type_cast_706_wire_constant <= "11001110";
    type_cast_708_wire_constant <= "11001111";
    type_cast_716_wire_constant <= "10110100";
    type_cast_718_wire_constant <= "11110000";
    type_cast_726_wire_constant <= "01110011";
    type_cast_728_wire_constant <= "11100110";
    type_cast_736_wire_constant <= "10101100";
    type_cast_738_wire_constant <= "10010110";
    type_cast_746_wire_constant <= "00100010";
    type_cast_748_wire_constant <= "01110100";
    type_cast_756_wire_constant <= "10101101";
    type_cast_758_wire_constant <= "11100111";
    type_cast_766_wire_constant <= "10000101";
    type_cast_768_wire_constant <= "00110101";
    type_cast_76_wire_constant <= "11110011";
    type_cast_776_wire_constant <= "11111001";
    type_cast_778_wire_constant <= "11100010";
    type_cast_786_wire_constant <= "11101000";
    type_cast_788_wire_constant <= "00110111";
    type_cast_78_wire_constant <= "10000001";
    type_cast_796_wire_constant <= "01110101";
    type_cast_798_wire_constant <= "00011100";
    type_cast_806_wire_constant <= "01101110";
    type_cast_808_wire_constant <= "11011111";
    type_cast_816_wire_constant <= "11110001";
    type_cast_818_wire_constant <= "01000111";
    type_cast_826_wire_constant <= "01110001";
    type_cast_828_wire_constant <= "00011010";
    type_cast_836_wire_constant <= "00101001";
    type_cast_838_wire_constant <= "00011101";
    type_cast_846_wire_constant <= "10001001";
    type_cast_848_wire_constant <= "11000101";
    type_cast_856_wire_constant <= "10110111";
    type_cast_858_wire_constant <= "01101111";
    type_cast_866_wire_constant <= "00001110";
    type_cast_868_wire_constant <= "01100010";
    type_cast_86_wire_constant <= "11111011";
    type_cast_876_wire_constant <= "00011000";
    type_cast_878_wire_constant <= "10101010";
    type_cast_886_wire_constant <= "00011011";
    type_cast_888_wire_constant <= "10111110";
    type_cast_88_wire_constant <= "11010111";
    type_cast_896_wire_constant <= "01010110";
    type_cast_898_wire_constant <= "11111100";
    type_cast_906_wire_constant <= "01001011";
    type_cast_908_wire_constant <= "00111110";
    type_cast_916_wire_constant <= "11010010";
    type_cast_918_wire_constant <= "11000110";
    type_cast_926_wire_constant <= "00100000";
    type_cast_928_wire_constant <= "01111001";
    type_cast_936_wire_constant <= "11011011";
    type_cast_938_wire_constant <= "10011010";
    type_cast_946_wire_constant <= "11111110";
    type_cast_948_wire_constant <= "11000000";
    type_cast_956_wire_constant <= "11001101";
    type_cast_958_wire_constant <= "01111000";
    type_cast_966_wire_constant <= "11110100";
    type_cast_968_wire_constant <= "01011010";
    type_cast_96_wire_constant <= "11100011";
    type_cast_976_wire_constant <= "11011101";
    type_cast_978_wire_constant <= "00011111";
    type_cast_986_wire_constant <= "00110011";
    type_cast_988_wire_constant <= "10101000";
    type_cast_98_wire_constant <= "01111100";
    type_cast_996_wire_constant <= "00000111";
    type_cast_998_wire_constant <= "10001000";
    -- logger for split-operator MUX_1009_inst flow-through 
    process(IMA99_1010) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1009_inst:flowthrough inputs: " & " BITSEL_u8_u1_1004_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1004_wire) & " type_cast_1006_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1006_wire_constant) & " type_cast_1008_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1008_wire_constant) & " outputs:" & " IMA99_1010= "  & Convert_SLV_To_Hex_String(IMA99_1010));
      --
    end process; 
    -- flow-through select operator MUX_1009_inst
    IMA99_1010 <= type_cast_1006_wire_constant when (BITSEL_u8_u1_1004_wire(0) /=  '0') else type_cast_1008_wire_constant;
    -- logger for split-operator MUX_1019_inst flow-through 
    process(IMA100_1020) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1019_inst:flowthrough inputs: " & " BITSEL_u8_u1_1014_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1014_wire) & " type_cast_1016_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1016_wire_constant) & " type_cast_1018_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1018_wire_constant) & " outputs:" & " IMA100_1020= "  & Convert_SLV_To_Hex_String(IMA100_1020));
      --
    end process; 
    -- flow-through select operator MUX_1019_inst
    IMA100_1020 <= type_cast_1016_wire_constant when (BITSEL_u8_u1_1014_wire(0) /=  '0') else type_cast_1018_wire_constant;
    -- logger for split-operator MUX_1029_inst flow-through 
    process(IMA101_1030) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1029_inst:flowthrough inputs: " & " BITSEL_u8_u1_1024_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1024_wire) & " type_cast_1026_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1026_wire_constant) & " type_cast_1028_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1028_wire_constant) & " outputs:" & " IMA101_1030= "  & Convert_SLV_To_Hex_String(IMA101_1030));
      --
    end process; 
    -- flow-through select operator MUX_1029_inst
    IMA101_1030 <= type_cast_1026_wire_constant when (BITSEL_u8_u1_1024_wire(0) /=  '0') else type_cast_1028_wire_constant;
    -- logger for split-operator MUX_1039_inst flow-through 
    process(IMA102_1040) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1039_inst:flowthrough inputs: " & " BITSEL_u8_u1_1034_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1034_wire) & " type_cast_1036_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1036_wire_constant) & " type_cast_1038_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1038_wire_constant) & " outputs:" & " IMA102_1040= "  & Convert_SLV_To_Hex_String(IMA102_1040));
      --
    end process; 
    -- flow-through select operator MUX_1039_inst
    IMA102_1040 <= type_cast_1036_wire_constant when (BITSEL_u8_u1_1034_wire(0) /=  '0') else type_cast_1038_wire_constant;
    -- logger for split-operator MUX_1049_inst flow-through 
    process(IMA103_1050) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1049_inst:flowthrough inputs: " & " BITSEL_u8_u1_1044_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1044_wire) & " type_cast_1046_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1046_wire_constant) & " type_cast_1048_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1048_wire_constant) & " outputs:" & " IMA103_1050= "  & Convert_SLV_To_Hex_String(IMA103_1050));
      --
    end process; 
    -- flow-through select operator MUX_1049_inst
    IMA103_1050 <= type_cast_1046_wire_constant when (BITSEL_u8_u1_1044_wire(0) /=  '0') else type_cast_1048_wire_constant;
    -- logger for split-operator MUX_1059_inst flow-through 
    process(IMA104_1060) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1059_inst:flowthrough inputs: " & " BITSEL_u8_u1_1054_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1054_wire) & " type_cast_1056_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1056_wire_constant) & " type_cast_1058_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1058_wire_constant) & " outputs:" & " IMA104_1060= "  & Convert_SLV_To_Hex_String(IMA104_1060));
      --
    end process; 
    -- flow-through select operator MUX_1059_inst
    IMA104_1060 <= type_cast_1056_wire_constant when (BITSEL_u8_u1_1054_wire(0) /=  '0') else type_cast_1058_wire_constant;
    -- logger for split-operator MUX_1069_inst flow-through 
    process(IMA105_1070) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1069_inst:flowthrough inputs: " & " BITSEL_u8_u1_1064_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1064_wire) & " type_cast_1066_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1066_wire_constant) & " type_cast_1068_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1068_wire_constant) & " outputs:" & " IMA105_1070= "  & Convert_SLV_To_Hex_String(IMA105_1070));
      --
    end process; 
    -- flow-through select operator MUX_1069_inst
    IMA105_1070 <= type_cast_1066_wire_constant when (BITSEL_u8_u1_1064_wire(0) /=  '0') else type_cast_1068_wire_constant;
    -- logger for split-operator MUX_1079_inst flow-through 
    process(IMA106_1080) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1079_inst:flowthrough inputs: " & " BITSEL_u8_u1_1074_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1074_wire) & " type_cast_1076_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1076_wire_constant) & " type_cast_1078_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1078_wire_constant) & " outputs:" & " IMA106_1080= "  & Convert_SLV_To_Hex_String(IMA106_1080));
      --
    end process; 
    -- flow-through select operator MUX_1079_inst
    IMA106_1080 <= type_cast_1076_wire_constant when (BITSEL_u8_u1_1074_wire(0) /=  '0') else type_cast_1078_wire_constant;
    -- logger for split-operator MUX_1089_inst flow-through 
    process(IMA107_1090) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1089_inst:flowthrough inputs: " & " BITSEL_u8_u1_1084_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1084_wire) & " type_cast_1086_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1086_wire_constant) & " type_cast_1088_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1088_wire_constant) & " outputs:" & " IMA107_1090= "  & Convert_SLV_To_Hex_String(IMA107_1090));
      --
    end process; 
    -- flow-through select operator MUX_1089_inst
    IMA107_1090 <= type_cast_1086_wire_constant when (BITSEL_u8_u1_1084_wire(0) /=  '0') else type_cast_1088_wire_constant;
    -- logger for split-operator MUX_1099_inst flow-through 
    process(IMA108_1100) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1099_inst:flowthrough inputs: " & " BITSEL_u8_u1_1094_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1094_wire) & " type_cast_1096_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1096_wire_constant) & " type_cast_1098_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1098_wire_constant) & " outputs:" & " IMA108_1100= "  & Convert_SLV_To_Hex_String(IMA108_1100));
      --
    end process; 
    -- flow-through select operator MUX_1099_inst
    IMA108_1100 <= type_cast_1096_wire_constant when (BITSEL_u8_u1_1094_wire(0) /=  '0') else type_cast_1098_wire_constant;
    -- logger for split-operator MUX_109_inst flow-through 
    process(IMA9_110) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_109_inst:flowthrough inputs: " & " BITSEL_u8_u1_104_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_104_wire) & " type_cast_106_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_106_wire_constant) & " type_cast_108_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_108_wire_constant) & " outputs:" & " IMA9_110= "  & Convert_SLV_To_Hex_String(IMA9_110));
      --
    end process; 
    -- flow-through select operator MUX_109_inst
    IMA9_110 <= type_cast_106_wire_constant when (BITSEL_u8_u1_104_wire(0) /=  '0') else type_cast_108_wire_constant;
    -- logger for split-operator MUX_1109_inst flow-through 
    process(IMA109_1110) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1109_inst:flowthrough inputs: " & " BITSEL_u8_u1_1104_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1104_wire) & " type_cast_1106_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1106_wire_constant) & " type_cast_1108_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1108_wire_constant) & " outputs:" & " IMA109_1110= "  & Convert_SLV_To_Hex_String(IMA109_1110));
      --
    end process; 
    -- flow-through select operator MUX_1109_inst
    IMA109_1110 <= type_cast_1106_wire_constant when (BITSEL_u8_u1_1104_wire(0) /=  '0') else type_cast_1108_wire_constant;
    -- logger for split-operator MUX_1119_inst flow-through 
    process(IMA110_1120) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1119_inst:flowthrough inputs: " & " BITSEL_u8_u1_1114_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1114_wire) & " type_cast_1116_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1116_wire_constant) & " type_cast_1118_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1118_wire_constant) & " outputs:" & " IMA110_1120= "  & Convert_SLV_To_Hex_String(IMA110_1120));
      --
    end process; 
    -- flow-through select operator MUX_1119_inst
    IMA110_1120 <= type_cast_1116_wire_constant when (BITSEL_u8_u1_1114_wire(0) /=  '0') else type_cast_1118_wire_constant;
    -- logger for split-operator MUX_1129_inst flow-through 
    process(IMA111_1130) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1129_inst:flowthrough inputs: " & " BITSEL_u8_u1_1124_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1124_wire) & " type_cast_1126_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1126_wire_constant) & " type_cast_1128_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1128_wire_constant) & " outputs:" & " IMA111_1130= "  & Convert_SLV_To_Hex_String(IMA111_1130));
      --
    end process; 
    -- flow-through select operator MUX_1129_inst
    IMA111_1130 <= type_cast_1126_wire_constant when (BITSEL_u8_u1_1124_wire(0) /=  '0') else type_cast_1128_wire_constant;
    -- logger for split-operator MUX_1139_inst flow-through 
    process(IMA112_1140) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1139_inst:flowthrough inputs: " & " BITSEL_u8_u1_1134_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1134_wire) & " type_cast_1136_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1136_wire_constant) & " type_cast_1138_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1138_wire_constant) & " outputs:" & " IMA112_1140= "  & Convert_SLV_To_Hex_String(IMA112_1140));
      --
    end process; 
    -- flow-through select operator MUX_1139_inst
    IMA112_1140 <= type_cast_1136_wire_constant when (BITSEL_u8_u1_1134_wire(0) /=  '0') else type_cast_1138_wire_constant;
    -- logger for split-operator MUX_1149_inst flow-through 
    process(IMA113_1150) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1149_inst:flowthrough inputs: " & " BITSEL_u8_u1_1144_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1144_wire) & " type_cast_1146_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1146_wire_constant) & " type_cast_1148_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1148_wire_constant) & " outputs:" & " IMA113_1150= "  & Convert_SLV_To_Hex_String(IMA113_1150));
      --
    end process; 
    -- flow-through select operator MUX_1149_inst
    IMA113_1150 <= type_cast_1146_wire_constant when (BITSEL_u8_u1_1144_wire(0) /=  '0') else type_cast_1148_wire_constant;
    -- logger for split-operator MUX_1159_inst flow-through 
    process(IMA114_1160) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1159_inst:flowthrough inputs: " & " BITSEL_u8_u1_1154_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1154_wire) & " type_cast_1156_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1156_wire_constant) & " type_cast_1158_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1158_wire_constant) & " outputs:" & " IMA114_1160= "  & Convert_SLV_To_Hex_String(IMA114_1160));
      --
    end process; 
    -- flow-through select operator MUX_1159_inst
    IMA114_1160 <= type_cast_1156_wire_constant when (BITSEL_u8_u1_1154_wire(0) /=  '0') else type_cast_1158_wire_constant;
    -- logger for split-operator MUX_1169_inst flow-through 
    process(IMA115_1170) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1169_inst:flowthrough inputs: " & " BITSEL_u8_u1_1164_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1164_wire) & " type_cast_1166_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1166_wire_constant) & " type_cast_1168_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1168_wire_constant) & " outputs:" & " IMA115_1170= "  & Convert_SLV_To_Hex_String(IMA115_1170));
      --
    end process; 
    -- flow-through select operator MUX_1169_inst
    IMA115_1170 <= type_cast_1166_wire_constant when (BITSEL_u8_u1_1164_wire(0) /=  '0') else type_cast_1168_wire_constant;
    -- logger for split-operator MUX_1179_inst flow-through 
    process(IMA116_1180) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1179_inst:flowthrough inputs: " & " BITSEL_u8_u1_1174_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1174_wire) & " type_cast_1176_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1176_wire_constant) & " type_cast_1178_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1178_wire_constant) & " outputs:" & " IMA116_1180= "  & Convert_SLV_To_Hex_String(IMA116_1180));
      --
    end process; 
    -- flow-through select operator MUX_1179_inst
    IMA116_1180 <= type_cast_1176_wire_constant when (BITSEL_u8_u1_1174_wire(0) /=  '0') else type_cast_1178_wire_constant;
    -- logger for split-operator MUX_1189_inst flow-through 
    process(IMA117_1190) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1189_inst:flowthrough inputs: " & " BITSEL_u8_u1_1184_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1184_wire) & " type_cast_1186_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1186_wire_constant) & " type_cast_1188_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1188_wire_constant) & " outputs:" & " IMA117_1190= "  & Convert_SLV_To_Hex_String(IMA117_1190));
      --
    end process; 
    -- flow-through select operator MUX_1189_inst
    IMA117_1190 <= type_cast_1186_wire_constant when (BITSEL_u8_u1_1184_wire(0) /=  '0') else type_cast_1188_wire_constant;
    -- logger for split-operator MUX_1199_inst flow-through 
    process(IMA118_1200) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1199_inst:flowthrough inputs: " & " BITSEL_u8_u1_1194_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1194_wire) & " type_cast_1196_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1196_wire_constant) & " type_cast_1198_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1198_wire_constant) & " outputs:" & " IMA118_1200= "  & Convert_SLV_To_Hex_String(IMA118_1200));
      --
    end process; 
    -- flow-through select operator MUX_1199_inst
    IMA118_1200 <= type_cast_1196_wire_constant when (BITSEL_u8_u1_1194_wire(0) /=  '0') else type_cast_1198_wire_constant;
    -- logger for split-operator MUX_119_inst flow-through 
    process(IMA10_120) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_119_inst:flowthrough inputs: " & " BITSEL_u8_u1_114_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_114_wire) & " type_cast_116_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_116_wire_constant) & " type_cast_118_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_118_wire_constant) & " outputs:" & " IMA10_120= "  & Convert_SLV_To_Hex_String(IMA10_120));
      --
    end process; 
    -- flow-through select operator MUX_119_inst
    IMA10_120 <= type_cast_116_wire_constant when (BITSEL_u8_u1_114_wire(0) /=  '0') else type_cast_118_wire_constant;
    -- logger for split-operator MUX_1209_inst flow-through 
    process(IMA119_1210) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1209_inst:flowthrough inputs: " & " BITSEL_u8_u1_1204_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1204_wire) & " type_cast_1206_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1206_wire_constant) & " type_cast_1208_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1208_wire_constant) & " outputs:" & " IMA119_1210= "  & Convert_SLV_To_Hex_String(IMA119_1210));
      --
    end process; 
    -- flow-through select operator MUX_1209_inst
    IMA119_1210 <= type_cast_1206_wire_constant when (BITSEL_u8_u1_1204_wire(0) /=  '0') else type_cast_1208_wire_constant;
    -- logger for split-operator MUX_1219_inst flow-through 
    process(IMA120_1220) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1219_inst:flowthrough inputs: " & " BITSEL_u8_u1_1214_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1214_wire) & " type_cast_1216_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1216_wire_constant) & " type_cast_1218_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1218_wire_constant) & " outputs:" & " IMA120_1220= "  & Convert_SLV_To_Hex_String(IMA120_1220));
      --
    end process; 
    -- flow-through select operator MUX_1219_inst
    IMA120_1220 <= type_cast_1216_wire_constant when (BITSEL_u8_u1_1214_wire(0) /=  '0') else type_cast_1218_wire_constant;
    -- logger for split-operator MUX_1229_inst flow-through 
    process(IMA121_1230) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1229_inst:flowthrough inputs: " & " BITSEL_u8_u1_1224_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1224_wire) & " type_cast_1226_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1226_wire_constant) & " type_cast_1228_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1228_wire_constant) & " outputs:" & " IMA121_1230= "  & Convert_SLV_To_Hex_String(IMA121_1230));
      --
    end process; 
    -- flow-through select operator MUX_1229_inst
    IMA121_1230 <= type_cast_1226_wire_constant when (BITSEL_u8_u1_1224_wire(0) /=  '0') else type_cast_1228_wire_constant;
    -- logger for split-operator MUX_1239_inst flow-through 
    process(IMA122_1240) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1239_inst:flowthrough inputs: " & " BITSEL_u8_u1_1234_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1234_wire) & " type_cast_1236_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1236_wire_constant) & " type_cast_1238_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1238_wire_constant) & " outputs:" & " IMA122_1240= "  & Convert_SLV_To_Hex_String(IMA122_1240));
      --
    end process; 
    -- flow-through select operator MUX_1239_inst
    IMA122_1240 <= type_cast_1236_wire_constant when (BITSEL_u8_u1_1234_wire(0) /=  '0') else type_cast_1238_wire_constant;
    -- logger for split-operator MUX_1249_inst flow-through 
    process(IMA123_1250) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1249_inst:flowthrough inputs: " & " BITSEL_u8_u1_1244_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1244_wire) & " type_cast_1246_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1246_wire_constant) & " type_cast_1248_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1248_wire_constant) & " outputs:" & " IMA123_1250= "  & Convert_SLV_To_Hex_String(IMA123_1250));
      --
    end process; 
    -- flow-through select operator MUX_1249_inst
    IMA123_1250 <= type_cast_1246_wire_constant when (BITSEL_u8_u1_1244_wire(0) /=  '0') else type_cast_1248_wire_constant;
    -- logger for split-operator MUX_1259_inst flow-through 
    process(IMA124_1260) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1259_inst:flowthrough inputs: " & " BITSEL_u8_u1_1254_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1254_wire) & " type_cast_1256_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1256_wire_constant) & " type_cast_1258_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1258_wire_constant) & " outputs:" & " IMA124_1260= "  & Convert_SLV_To_Hex_String(IMA124_1260));
      --
    end process; 
    -- flow-through select operator MUX_1259_inst
    IMA124_1260 <= type_cast_1256_wire_constant when (BITSEL_u8_u1_1254_wire(0) /=  '0') else type_cast_1258_wire_constant;
    -- logger for split-operator MUX_1269_inst flow-through 
    process(IMA125_1270) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1269_inst:flowthrough inputs: " & " BITSEL_u8_u1_1264_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1264_wire) & " type_cast_1266_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1266_wire_constant) & " type_cast_1268_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1268_wire_constant) & " outputs:" & " IMA125_1270= "  & Convert_SLV_To_Hex_String(IMA125_1270));
      --
    end process; 
    -- flow-through select operator MUX_1269_inst
    IMA125_1270 <= type_cast_1266_wire_constant when (BITSEL_u8_u1_1264_wire(0) /=  '0') else type_cast_1268_wire_constant;
    -- logger for split-operator MUX_1279_inst flow-through 
    process(IMA126_1280) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1279_inst:flowthrough inputs: " & " BITSEL_u8_u1_1274_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1274_wire) & " type_cast_1276_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1276_wire_constant) & " type_cast_1278_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1278_wire_constant) & " outputs:" & " IMA126_1280= "  & Convert_SLV_To_Hex_String(IMA126_1280));
      --
    end process; 
    -- flow-through select operator MUX_1279_inst
    IMA126_1280 <= type_cast_1276_wire_constant when (BITSEL_u8_u1_1274_wire(0) /=  '0') else type_cast_1278_wire_constant;
    -- logger for split-operator MUX_1289_inst flow-through 
    process(IMA127_1290) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1289_inst:flowthrough inputs: " & " BITSEL_u8_u1_1284_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1284_wire) & " type_cast_1286_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1286_wire_constant) & " type_cast_1288_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1288_wire_constant) & " outputs:" & " IMA127_1290= "  & Convert_SLV_To_Hex_String(IMA127_1290));
      --
    end process; 
    -- flow-through select operator MUX_1289_inst
    IMA127_1290 <= type_cast_1286_wire_constant when (BITSEL_u8_u1_1284_wire(0) /=  '0') else type_cast_1288_wire_constant;
    -- logger for split-operator MUX_1297_inst flow-through 
    process(IMB0_1298) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1297_inst:flowthrough inputs: " & " BITSEL_u8_u1_1294_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1294_wire) & " IMA1_30 = "& Convert_SLV_To_Hex_String(IMA1_30) & " IMA0_20 = "& Convert_SLV_To_Hex_String(IMA0_20) & " outputs:" & " IMB0_1298= "  & Convert_SLV_To_Hex_String(IMB0_1298));
      --
    end process; 
    -- flow-through select operator MUX_1297_inst
    IMB0_1298 <= IMA1_30 when (BITSEL_u8_u1_1294_wire(0) /=  '0') else IMA0_20;
    -- logger for split-operator MUX_129_inst flow-through 
    process(IMA11_130) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_129_inst:flowthrough inputs: " & " BITSEL_u8_u1_124_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_124_wire) & " type_cast_126_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_126_wire_constant) & " type_cast_128_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_128_wire_constant) & " outputs:" & " IMA11_130= "  & Convert_SLV_To_Hex_String(IMA11_130));
      --
    end process; 
    -- flow-through select operator MUX_129_inst
    IMA11_130 <= type_cast_126_wire_constant when (BITSEL_u8_u1_124_wire(0) /=  '0') else type_cast_128_wire_constant;
    -- logger for split-operator MUX_1305_inst flow-through 
    process(IMB1_1306) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1305_inst:flowthrough inputs: " & " BITSEL_u8_u1_1302_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1302_wire) & " IMA3_50 = "& Convert_SLV_To_Hex_String(IMA3_50) & " IMA2_40 = "& Convert_SLV_To_Hex_String(IMA2_40) & " outputs:" & " IMB1_1306= "  & Convert_SLV_To_Hex_String(IMB1_1306));
      --
    end process; 
    -- flow-through select operator MUX_1305_inst
    IMB1_1306 <= IMA3_50 when (BITSEL_u8_u1_1302_wire(0) /=  '0') else IMA2_40;
    -- logger for split-operator MUX_1313_inst flow-through 
    process(IMB2_1314) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1313_inst:flowthrough inputs: " & " BITSEL_u8_u1_1310_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1310_wire) & " IMA5_70 = "& Convert_SLV_To_Hex_String(IMA5_70) & " IMA4_60 = "& Convert_SLV_To_Hex_String(IMA4_60) & " outputs:" & " IMB2_1314= "  & Convert_SLV_To_Hex_String(IMB2_1314));
      --
    end process; 
    -- flow-through select operator MUX_1313_inst
    IMB2_1314 <= IMA5_70 when (BITSEL_u8_u1_1310_wire(0) /=  '0') else IMA4_60;
    -- logger for split-operator MUX_1321_inst flow-through 
    process(IMB3_1322) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1321_inst:flowthrough inputs: " & " BITSEL_u8_u1_1318_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1318_wire) & " IMA7_90 = "& Convert_SLV_To_Hex_String(IMA7_90) & " IMA6_80 = "& Convert_SLV_To_Hex_String(IMA6_80) & " outputs:" & " IMB3_1322= "  & Convert_SLV_To_Hex_String(IMB3_1322));
      --
    end process; 
    -- flow-through select operator MUX_1321_inst
    IMB3_1322 <= IMA7_90 when (BITSEL_u8_u1_1318_wire(0) /=  '0') else IMA6_80;
    -- logger for split-operator MUX_1329_inst flow-through 
    process(IMB4_1330) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1329_inst:flowthrough inputs: " & " BITSEL_u8_u1_1326_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1326_wire) & " IMA9_110 = "& Convert_SLV_To_Hex_String(IMA9_110) & " IMA8_100 = "& Convert_SLV_To_Hex_String(IMA8_100) & " outputs:" & " IMB4_1330= "  & Convert_SLV_To_Hex_String(IMB4_1330));
      --
    end process; 
    -- flow-through select operator MUX_1329_inst
    IMB4_1330 <= IMA9_110 when (BITSEL_u8_u1_1326_wire(0) /=  '0') else IMA8_100;
    -- logger for split-operator MUX_1337_inst flow-through 
    process(IMB5_1338) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1337_inst:flowthrough inputs: " & " BITSEL_u8_u1_1334_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1334_wire) & " IMA11_130 = "& Convert_SLV_To_Hex_String(IMA11_130) & " IMA10_120 = "& Convert_SLV_To_Hex_String(IMA10_120) & " outputs:" & " IMB5_1338= "  & Convert_SLV_To_Hex_String(IMB5_1338));
      --
    end process; 
    -- flow-through select operator MUX_1337_inst
    IMB5_1338 <= IMA11_130 when (BITSEL_u8_u1_1334_wire(0) /=  '0') else IMA10_120;
    -- logger for split-operator MUX_1345_inst flow-through 
    process(IMB6_1346) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1345_inst:flowthrough inputs: " & " BITSEL_u8_u1_1342_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1342_wire) & " IMA13_150 = "& Convert_SLV_To_Hex_String(IMA13_150) & " IMA12_140 = "& Convert_SLV_To_Hex_String(IMA12_140) & " outputs:" & " IMB6_1346= "  & Convert_SLV_To_Hex_String(IMB6_1346));
      --
    end process; 
    -- flow-through select operator MUX_1345_inst
    IMB6_1346 <= IMA13_150 when (BITSEL_u8_u1_1342_wire(0) /=  '0') else IMA12_140;
    -- logger for split-operator MUX_1353_inst flow-through 
    process(IMB7_1354) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1353_inst:flowthrough inputs: " & " BITSEL_u8_u1_1350_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1350_wire) & " IMA15_170 = "& Convert_SLV_To_Hex_String(IMA15_170) & " IMA14_160 = "& Convert_SLV_To_Hex_String(IMA14_160) & " outputs:" & " IMB7_1354= "  & Convert_SLV_To_Hex_String(IMB7_1354));
      --
    end process; 
    -- flow-through select operator MUX_1353_inst
    IMB7_1354 <= IMA15_170 when (BITSEL_u8_u1_1350_wire(0) /=  '0') else IMA14_160;
    -- logger for split-operator MUX_1361_inst flow-through 
    process(IMB8_1362) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1361_inst:flowthrough inputs: " & " BITSEL_u8_u1_1358_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1358_wire) & " IMA17_190 = "& Convert_SLV_To_Hex_String(IMA17_190) & " IMA16_180 = "& Convert_SLV_To_Hex_String(IMA16_180) & " outputs:" & " IMB8_1362= "  & Convert_SLV_To_Hex_String(IMB8_1362));
      --
    end process; 
    -- flow-through select operator MUX_1361_inst
    IMB8_1362 <= IMA17_190 when (BITSEL_u8_u1_1358_wire(0) /=  '0') else IMA16_180;
    -- logger for split-operator MUX_1369_inst flow-through 
    process(IMB9_1370) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1369_inst:flowthrough inputs: " & " BITSEL_u8_u1_1366_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1366_wire) & " IMA19_210 = "& Convert_SLV_To_Hex_String(IMA19_210) & " IMA18_200 = "& Convert_SLV_To_Hex_String(IMA18_200) & " outputs:" & " IMB9_1370= "  & Convert_SLV_To_Hex_String(IMB9_1370));
      --
    end process; 
    -- flow-through select operator MUX_1369_inst
    IMB9_1370 <= IMA19_210 when (BITSEL_u8_u1_1366_wire(0) /=  '0') else IMA18_200;
    -- logger for split-operator MUX_1377_inst flow-through 
    process(IMB10_1378) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1377_inst:flowthrough inputs: " & " BITSEL_u8_u1_1374_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1374_wire) & " IMA21_230 = "& Convert_SLV_To_Hex_String(IMA21_230) & " IMA20_220 = "& Convert_SLV_To_Hex_String(IMA20_220) & " outputs:" & " IMB10_1378= "  & Convert_SLV_To_Hex_String(IMB10_1378));
      --
    end process; 
    -- flow-through select operator MUX_1377_inst
    IMB10_1378 <= IMA21_230 when (BITSEL_u8_u1_1374_wire(0) /=  '0') else IMA20_220;
    -- logger for split-operator MUX_1385_inst flow-through 
    process(IMB11_1386) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1385_inst:flowthrough inputs: " & " BITSEL_u8_u1_1382_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1382_wire) & " IMA23_250 = "& Convert_SLV_To_Hex_String(IMA23_250) & " IMA22_240 = "& Convert_SLV_To_Hex_String(IMA22_240) & " outputs:" & " IMB11_1386= "  & Convert_SLV_To_Hex_String(IMB11_1386));
      --
    end process; 
    -- flow-through select operator MUX_1385_inst
    IMB11_1386 <= IMA23_250 when (BITSEL_u8_u1_1382_wire(0) /=  '0') else IMA22_240;
    -- logger for split-operator MUX_1393_inst flow-through 
    process(IMB12_1394) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1393_inst:flowthrough inputs: " & " BITSEL_u8_u1_1390_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1390_wire) & " IMA25_270 = "& Convert_SLV_To_Hex_String(IMA25_270) & " IMA24_260 = "& Convert_SLV_To_Hex_String(IMA24_260) & " outputs:" & " IMB12_1394= "  & Convert_SLV_To_Hex_String(IMB12_1394));
      --
    end process; 
    -- flow-through select operator MUX_1393_inst
    IMB12_1394 <= IMA25_270 when (BITSEL_u8_u1_1390_wire(0) /=  '0') else IMA24_260;
    -- logger for split-operator MUX_139_inst flow-through 
    process(IMA12_140) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_139_inst:flowthrough inputs: " & " BITSEL_u8_u1_134_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_134_wire) & " type_cast_136_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_136_wire_constant) & " type_cast_138_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_138_wire_constant) & " outputs:" & " IMA12_140= "  & Convert_SLV_To_Hex_String(IMA12_140));
      --
    end process; 
    -- flow-through select operator MUX_139_inst
    IMA12_140 <= type_cast_136_wire_constant when (BITSEL_u8_u1_134_wire(0) /=  '0') else type_cast_138_wire_constant;
    -- logger for split-operator MUX_1401_inst flow-through 
    process(IMB13_1402) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1401_inst:flowthrough inputs: " & " BITSEL_u8_u1_1398_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1398_wire) & " IMA27_290 = "& Convert_SLV_To_Hex_String(IMA27_290) & " IMA26_280 = "& Convert_SLV_To_Hex_String(IMA26_280) & " outputs:" & " IMB13_1402= "  & Convert_SLV_To_Hex_String(IMB13_1402));
      --
    end process; 
    -- flow-through select operator MUX_1401_inst
    IMB13_1402 <= IMA27_290 when (BITSEL_u8_u1_1398_wire(0) /=  '0') else IMA26_280;
    -- logger for split-operator MUX_1409_inst flow-through 
    process(IMB14_1410) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1409_inst:flowthrough inputs: " & " BITSEL_u8_u1_1406_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1406_wire) & " IMA29_310 = "& Convert_SLV_To_Hex_String(IMA29_310) & " IMA28_300 = "& Convert_SLV_To_Hex_String(IMA28_300) & " outputs:" & " IMB14_1410= "  & Convert_SLV_To_Hex_String(IMB14_1410));
      --
    end process; 
    -- flow-through select operator MUX_1409_inst
    IMB14_1410 <= IMA29_310 when (BITSEL_u8_u1_1406_wire(0) /=  '0') else IMA28_300;
    -- logger for split-operator MUX_1417_inst flow-through 
    process(IMB15_1418) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1417_inst:flowthrough inputs: " & " BITSEL_u8_u1_1414_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1414_wire) & " IMA31_330 = "& Convert_SLV_To_Hex_String(IMA31_330) & " IMA30_320 = "& Convert_SLV_To_Hex_String(IMA30_320) & " outputs:" & " IMB15_1418= "  & Convert_SLV_To_Hex_String(IMB15_1418));
      --
    end process; 
    -- flow-through select operator MUX_1417_inst
    IMB15_1418 <= IMA31_330 when (BITSEL_u8_u1_1414_wire(0) /=  '0') else IMA30_320;
    -- logger for split-operator MUX_1425_inst flow-through 
    process(IMB16_1426) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1425_inst:flowthrough inputs: " & " BITSEL_u8_u1_1422_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1422_wire) & " IMA33_350 = "& Convert_SLV_To_Hex_String(IMA33_350) & " IMA32_340 = "& Convert_SLV_To_Hex_String(IMA32_340) & " outputs:" & " IMB16_1426= "  & Convert_SLV_To_Hex_String(IMB16_1426));
      --
    end process; 
    -- flow-through select operator MUX_1425_inst
    IMB16_1426 <= IMA33_350 when (BITSEL_u8_u1_1422_wire(0) /=  '0') else IMA32_340;
    -- logger for split-operator MUX_1433_inst flow-through 
    process(IMB17_1434) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1433_inst:flowthrough inputs: " & " BITSEL_u8_u1_1430_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1430_wire) & " IMA35_370 = "& Convert_SLV_To_Hex_String(IMA35_370) & " IMA34_360 = "& Convert_SLV_To_Hex_String(IMA34_360) & " outputs:" & " IMB17_1434= "  & Convert_SLV_To_Hex_String(IMB17_1434));
      --
    end process; 
    -- flow-through select operator MUX_1433_inst
    IMB17_1434 <= IMA35_370 when (BITSEL_u8_u1_1430_wire(0) /=  '0') else IMA34_360;
    -- logger for split-operator MUX_1441_inst flow-through 
    process(IMB18_1442) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1441_inst:flowthrough inputs: " & " BITSEL_u8_u1_1438_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1438_wire) & " IMA37_390 = "& Convert_SLV_To_Hex_String(IMA37_390) & " IMA36_380 = "& Convert_SLV_To_Hex_String(IMA36_380) & " outputs:" & " IMB18_1442= "  & Convert_SLV_To_Hex_String(IMB18_1442));
      --
    end process; 
    -- flow-through select operator MUX_1441_inst
    IMB18_1442 <= IMA37_390 when (BITSEL_u8_u1_1438_wire(0) /=  '0') else IMA36_380;
    -- logger for split-operator MUX_1449_inst flow-through 
    process(IMB19_1450) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1449_inst:flowthrough inputs: " & " BITSEL_u8_u1_1446_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1446_wire) & " IMA39_410 = "& Convert_SLV_To_Hex_String(IMA39_410) & " IMA38_400 = "& Convert_SLV_To_Hex_String(IMA38_400) & " outputs:" & " IMB19_1450= "  & Convert_SLV_To_Hex_String(IMB19_1450));
      --
    end process; 
    -- flow-through select operator MUX_1449_inst
    IMB19_1450 <= IMA39_410 when (BITSEL_u8_u1_1446_wire(0) /=  '0') else IMA38_400;
    -- logger for split-operator MUX_1457_inst flow-through 
    process(IMB20_1458) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1457_inst:flowthrough inputs: " & " BITSEL_u8_u1_1454_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1454_wire) & " IMA41_430 = "& Convert_SLV_To_Hex_String(IMA41_430) & " IMA40_420 = "& Convert_SLV_To_Hex_String(IMA40_420) & " outputs:" & " IMB20_1458= "  & Convert_SLV_To_Hex_String(IMB20_1458));
      --
    end process; 
    -- flow-through select operator MUX_1457_inst
    IMB20_1458 <= IMA41_430 when (BITSEL_u8_u1_1454_wire(0) /=  '0') else IMA40_420;
    -- logger for split-operator MUX_1465_inst flow-through 
    process(IMB21_1466) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1465_inst:flowthrough inputs: " & " BITSEL_u8_u1_1462_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1462_wire) & " IMA43_450 = "& Convert_SLV_To_Hex_String(IMA43_450) & " IMA42_440 = "& Convert_SLV_To_Hex_String(IMA42_440) & " outputs:" & " IMB21_1466= "  & Convert_SLV_To_Hex_String(IMB21_1466));
      --
    end process; 
    -- flow-through select operator MUX_1465_inst
    IMB21_1466 <= IMA43_450 when (BITSEL_u8_u1_1462_wire(0) /=  '0') else IMA42_440;
    -- logger for split-operator MUX_1473_inst flow-through 
    process(IMB22_1474) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1473_inst:flowthrough inputs: " & " BITSEL_u8_u1_1470_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1470_wire) & " IMA45_470 = "& Convert_SLV_To_Hex_String(IMA45_470) & " IMA44_460 = "& Convert_SLV_To_Hex_String(IMA44_460) & " outputs:" & " IMB22_1474= "  & Convert_SLV_To_Hex_String(IMB22_1474));
      --
    end process; 
    -- flow-through select operator MUX_1473_inst
    IMB22_1474 <= IMA45_470 when (BITSEL_u8_u1_1470_wire(0) /=  '0') else IMA44_460;
    -- logger for split-operator MUX_1481_inst flow-through 
    process(IMB23_1482) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1481_inst:flowthrough inputs: " & " BITSEL_u8_u1_1478_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1478_wire) & " IMA47_490 = "& Convert_SLV_To_Hex_String(IMA47_490) & " IMA46_480 = "& Convert_SLV_To_Hex_String(IMA46_480) & " outputs:" & " IMB23_1482= "  & Convert_SLV_To_Hex_String(IMB23_1482));
      --
    end process; 
    -- flow-through select operator MUX_1481_inst
    IMB23_1482 <= IMA47_490 when (BITSEL_u8_u1_1478_wire(0) /=  '0') else IMA46_480;
    -- logger for split-operator MUX_1489_inst flow-through 
    process(IMB24_1490) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1489_inst:flowthrough inputs: " & " BITSEL_u8_u1_1486_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1486_wire) & " IMA49_510 = "& Convert_SLV_To_Hex_String(IMA49_510) & " IMA48_500 = "& Convert_SLV_To_Hex_String(IMA48_500) & " outputs:" & " IMB24_1490= "  & Convert_SLV_To_Hex_String(IMB24_1490));
      --
    end process; 
    -- flow-through select operator MUX_1489_inst
    IMB24_1490 <= IMA49_510 when (BITSEL_u8_u1_1486_wire(0) /=  '0') else IMA48_500;
    -- logger for split-operator MUX_1497_inst flow-through 
    process(IMB25_1498) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1497_inst:flowthrough inputs: " & " BITSEL_u8_u1_1494_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1494_wire) & " IMA51_530 = "& Convert_SLV_To_Hex_String(IMA51_530) & " IMA50_520 = "& Convert_SLV_To_Hex_String(IMA50_520) & " outputs:" & " IMB25_1498= "  & Convert_SLV_To_Hex_String(IMB25_1498));
      --
    end process; 
    -- flow-through select operator MUX_1497_inst
    IMB25_1498 <= IMA51_530 when (BITSEL_u8_u1_1494_wire(0) /=  '0') else IMA50_520;
    -- logger for split-operator MUX_149_inst flow-through 
    process(IMA13_150) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_149_inst:flowthrough inputs: " & " BITSEL_u8_u1_144_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_144_wire) & " type_cast_146_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_146_wire_constant) & " type_cast_148_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_148_wire_constant) & " outputs:" & " IMA13_150= "  & Convert_SLV_To_Hex_String(IMA13_150));
      --
    end process; 
    -- flow-through select operator MUX_149_inst
    IMA13_150 <= type_cast_146_wire_constant when (BITSEL_u8_u1_144_wire(0) /=  '0') else type_cast_148_wire_constant;
    -- logger for split-operator MUX_1505_inst flow-through 
    process(IMB26_1506) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1505_inst:flowthrough inputs: " & " BITSEL_u8_u1_1502_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1502_wire) & " IMA53_550 = "& Convert_SLV_To_Hex_String(IMA53_550) & " IMA52_540 = "& Convert_SLV_To_Hex_String(IMA52_540) & " outputs:" & " IMB26_1506= "  & Convert_SLV_To_Hex_String(IMB26_1506));
      --
    end process; 
    -- flow-through select operator MUX_1505_inst
    IMB26_1506 <= IMA53_550 when (BITSEL_u8_u1_1502_wire(0) /=  '0') else IMA52_540;
    -- logger for split-operator MUX_1513_inst flow-through 
    process(IMB27_1514) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1513_inst:flowthrough inputs: " & " BITSEL_u8_u1_1510_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1510_wire) & " IMA55_570 = "& Convert_SLV_To_Hex_String(IMA55_570) & " IMA54_560 = "& Convert_SLV_To_Hex_String(IMA54_560) & " outputs:" & " IMB27_1514= "  & Convert_SLV_To_Hex_String(IMB27_1514));
      --
    end process; 
    -- flow-through select operator MUX_1513_inst
    IMB27_1514 <= IMA55_570 when (BITSEL_u8_u1_1510_wire(0) /=  '0') else IMA54_560;
    -- logger for split-operator MUX_1521_inst flow-through 
    process(IMB28_1522) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1521_inst:flowthrough inputs: " & " BITSEL_u8_u1_1518_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1518_wire) & " IMA57_590 = "& Convert_SLV_To_Hex_String(IMA57_590) & " IMA56_580 = "& Convert_SLV_To_Hex_String(IMA56_580) & " outputs:" & " IMB28_1522= "  & Convert_SLV_To_Hex_String(IMB28_1522));
      --
    end process; 
    -- flow-through select operator MUX_1521_inst
    IMB28_1522 <= IMA57_590 when (BITSEL_u8_u1_1518_wire(0) /=  '0') else IMA56_580;
    -- logger for split-operator MUX_1529_inst flow-through 
    process(IMB29_1530) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1529_inst:flowthrough inputs: " & " BITSEL_u8_u1_1526_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1526_wire) & " IMA59_610 = "& Convert_SLV_To_Hex_String(IMA59_610) & " IMA58_600 = "& Convert_SLV_To_Hex_String(IMA58_600) & " outputs:" & " IMB29_1530= "  & Convert_SLV_To_Hex_String(IMB29_1530));
      --
    end process; 
    -- flow-through select operator MUX_1529_inst
    IMB29_1530 <= IMA59_610 when (BITSEL_u8_u1_1526_wire(0) /=  '0') else IMA58_600;
    -- logger for split-operator MUX_1537_inst flow-through 
    process(IMB30_1538) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1537_inst:flowthrough inputs: " & " BITSEL_u8_u1_1534_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1534_wire) & " IMA61_630 = "& Convert_SLV_To_Hex_String(IMA61_630) & " IMA60_620 = "& Convert_SLV_To_Hex_String(IMA60_620) & " outputs:" & " IMB30_1538= "  & Convert_SLV_To_Hex_String(IMB30_1538));
      --
    end process; 
    -- flow-through select operator MUX_1537_inst
    IMB30_1538 <= IMA61_630 when (BITSEL_u8_u1_1534_wire(0) /=  '0') else IMA60_620;
    -- logger for split-operator MUX_1545_inst flow-through 
    process(IMB31_1546) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1545_inst:flowthrough inputs: " & " BITSEL_u8_u1_1542_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1542_wire) & " IMA63_650 = "& Convert_SLV_To_Hex_String(IMA63_650) & " IMA62_640 = "& Convert_SLV_To_Hex_String(IMA62_640) & " outputs:" & " IMB31_1546= "  & Convert_SLV_To_Hex_String(IMB31_1546));
      --
    end process; 
    -- flow-through select operator MUX_1545_inst
    IMB31_1546 <= IMA63_650 when (BITSEL_u8_u1_1542_wire(0) /=  '0') else IMA62_640;
    -- logger for split-operator MUX_1553_inst flow-through 
    process(IMB32_1554) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1553_inst:flowthrough inputs: " & " BITSEL_u8_u1_1550_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1550_wire) & " IMA65_670 = "& Convert_SLV_To_Hex_String(IMA65_670) & " IMA64_660 = "& Convert_SLV_To_Hex_String(IMA64_660) & " outputs:" & " IMB32_1554= "  & Convert_SLV_To_Hex_String(IMB32_1554));
      --
    end process; 
    -- flow-through select operator MUX_1553_inst
    IMB32_1554 <= IMA65_670 when (BITSEL_u8_u1_1550_wire(0) /=  '0') else IMA64_660;
    -- logger for split-operator MUX_1561_inst flow-through 
    process(IMB33_1562) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1561_inst:flowthrough inputs: " & " BITSEL_u8_u1_1558_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1558_wire) & " IMA67_690 = "& Convert_SLV_To_Hex_String(IMA67_690) & " IMA66_680 = "& Convert_SLV_To_Hex_String(IMA66_680) & " outputs:" & " IMB33_1562= "  & Convert_SLV_To_Hex_String(IMB33_1562));
      --
    end process; 
    -- flow-through select operator MUX_1561_inst
    IMB33_1562 <= IMA67_690 when (BITSEL_u8_u1_1558_wire(0) /=  '0') else IMA66_680;
    -- logger for split-operator MUX_1569_inst flow-through 
    process(IMB34_1570) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1569_inst:flowthrough inputs: " & " BITSEL_u8_u1_1566_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1566_wire) & " IMA69_710 = "& Convert_SLV_To_Hex_String(IMA69_710) & " IMA68_700 = "& Convert_SLV_To_Hex_String(IMA68_700) & " outputs:" & " IMB34_1570= "  & Convert_SLV_To_Hex_String(IMB34_1570));
      --
    end process; 
    -- flow-through select operator MUX_1569_inst
    IMB34_1570 <= IMA69_710 when (BITSEL_u8_u1_1566_wire(0) /=  '0') else IMA68_700;
    -- logger for split-operator MUX_1577_inst flow-through 
    process(IMB35_1578) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1577_inst:flowthrough inputs: " & " BITSEL_u8_u1_1574_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1574_wire) & " IMA71_730 = "& Convert_SLV_To_Hex_String(IMA71_730) & " IMA70_720 = "& Convert_SLV_To_Hex_String(IMA70_720) & " outputs:" & " IMB35_1578= "  & Convert_SLV_To_Hex_String(IMB35_1578));
      --
    end process; 
    -- flow-through select operator MUX_1577_inst
    IMB35_1578 <= IMA71_730 when (BITSEL_u8_u1_1574_wire(0) /=  '0') else IMA70_720;
    -- logger for split-operator MUX_1585_inst flow-through 
    process(IMB36_1586) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1585_inst:flowthrough inputs: " & " BITSEL_u8_u1_1582_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1582_wire) & " IMA73_750 = "& Convert_SLV_To_Hex_String(IMA73_750) & " IMA72_740 = "& Convert_SLV_To_Hex_String(IMA72_740) & " outputs:" & " IMB36_1586= "  & Convert_SLV_To_Hex_String(IMB36_1586));
      --
    end process; 
    -- flow-through select operator MUX_1585_inst
    IMB36_1586 <= IMA73_750 when (BITSEL_u8_u1_1582_wire(0) /=  '0') else IMA72_740;
    -- logger for split-operator MUX_1593_inst flow-through 
    process(IMB37_1594) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1593_inst:flowthrough inputs: " & " BITSEL_u8_u1_1590_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1590_wire) & " IMA75_770 = "& Convert_SLV_To_Hex_String(IMA75_770) & " IMA74_760 = "& Convert_SLV_To_Hex_String(IMA74_760) & " outputs:" & " IMB37_1594= "  & Convert_SLV_To_Hex_String(IMB37_1594));
      --
    end process; 
    -- flow-through select operator MUX_1593_inst
    IMB37_1594 <= IMA75_770 when (BITSEL_u8_u1_1590_wire(0) /=  '0') else IMA74_760;
    -- logger for split-operator MUX_159_inst flow-through 
    process(IMA14_160) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_159_inst:flowthrough inputs: " & " BITSEL_u8_u1_154_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_154_wire) & " type_cast_156_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_156_wire_constant) & " type_cast_158_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_158_wire_constant) & " outputs:" & " IMA14_160= "  & Convert_SLV_To_Hex_String(IMA14_160));
      --
    end process; 
    -- flow-through select operator MUX_159_inst
    IMA14_160 <= type_cast_156_wire_constant when (BITSEL_u8_u1_154_wire(0) /=  '0') else type_cast_158_wire_constant;
    -- logger for split-operator MUX_1601_inst flow-through 
    process(IMB38_1602) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1601_inst:flowthrough inputs: " & " BITSEL_u8_u1_1598_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1598_wire) & " IMA77_790 = "& Convert_SLV_To_Hex_String(IMA77_790) & " IMA76_780 = "& Convert_SLV_To_Hex_String(IMA76_780) & " outputs:" & " IMB38_1602= "  & Convert_SLV_To_Hex_String(IMB38_1602));
      --
    end process; 
    -- flow-through select operator MUX_1601_inst
    IMB38_1602 <= IMA77_790 when (BITSEL_u8_u1_1598_wire(0) /=  '0') else IMA76_780;
    -- logger for split-operator MUX_1609_inst flow-through 
    process(IMB39_1610) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1609_inst:flowthrough inputs: " & " BITSEL_u8_u1_1606_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1606_wire) & " IMA79_810 = "& Convert_SLV_To_Hex_String(IMA79_810) & " IMA78_800 = "& Convert_SLV_To_Hex_String(IMA78_800) & " outputs:" & " IMB39_1610= "  & Convert_SLV_To_Hex_String(IMB39_1610));
      --
    end process; 
    -- flow-through select operator MUX_1609_inst
    IMB39_1610 <= IMA79_810 when (BITSEL_u8_u1_1606_wire(0) /=  '0') else IMA78_800;
    -- logger for split-operator MUX_1617_inst flow-through 
    process(IMB40_1618) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1617_inst:flowthrough inputs: " & " BITSEL_u8_u1_1614_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1614_wire) & " IMA81_830 = "& Convert_SLV_To_Hex_String(IMA81_830) & " IMA80_820 = "& Convert_SLV_To_Hex_String(IMA80_820) & " outputs:" & " IMB40_1618= "  & Convert_SLV_To_Hex_String(IMB40_1618));
      --
    end process; 
    -- flow-through select operator MUX_1617_inst
    IMB40_1618 <= IMA81_830 when (BITSEL_u8_u1_1614_wire(0) /=  '0') else IMA80_820;
    -- logger for split-operator MUX_1625_inst flow-through 
    process(IMB41_1626) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1625_inst:flowthrough inputs: " & " BITSEL_u8_u1_1622_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1622_wire) & " IMA83_850 = "& Convert_SLV_To_Hex_String(IMA83_850) & " IMA82_840 = "& Convert_SLV_To_Hex_String(IMA82_840) & " outputs:" & " IMB41_1626= "  & Convert_SLV_To_Hex_String(IMB41_1626));
      --
    end process; 
    -- flow-through select operator MUX_1625_inst
    IMB41_1626 <= IMA83_850 when (BITSEL_u8_u1_1622_wire(0) /=  '0') else IMA82_840;
    -- logger for split-operator MUX_1633_inst flow-through 
    process(IMB42_1634) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1633_inst:flowthrough inputs: " & " BITSEL_u8_u1_1630_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1630_wire) & " IMA85_870 = "& Convert_SLV_To_Hex_String(IMA85_870) & " IMA84_860 = "& Convert_SLV_To_Hex_String(IMA84_860) & " outputs:" & " IMB42_1634= "  & Convert_SLV_To_Hex_String(IMB42_1634));
      --
    end process; 
    -- flow-through select operator MUX_1633_inst
    IMB42_1634 <= IMA85_870 when (BITSEL_u8_u1_1630_wire(0) /=  '0') else IMA84_860;
    -- logger for split-operator MUX_1641_inst flow-through 
    process(IMB43_1642) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1641_inst:flowthrough inputs: " & " BITSEL_u8_u1_1638_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1638_wire) & " IMA87_890 = "& Convert_SLV_To_Hex_String(IMA87_890) & " IMA86_880 = "& Convert_SLV_To_Hex_String(IMA86_880) & " outputs:" & " IMB43_1642= "  & Convert_SLV_To_Hex_String(IMB43_1642));
      --
    end process; 
    -- flow-through select operator MUX_1641_inst
    IMB43_1642 <= IMA87_890 when (BITSEL_u8_u1_1638_wire(0) /=  '0') else IMA86_880;
    -- logger for split-operator MUX_1649_inst flow-through 
    process(IMB44_1650) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1649_inst:flowthrough inputs: " & " BITSEL_u8_u1_1646_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1646_wire) & " IMA89_910 = "& Convert_SLV_To_Hex_String(IMA89_910) & " IMA88_900 = "& Convert_SLV_To_Hex_String(IMA88_900) & " outputs:" & " IMB44_1650= "  & Convert_SLV_To_Hex_String(IMB44_1650));
      --
    end process; 
    -- flow-through select operator MUX_1649_inst
    IMB44_1650 <= IMA89_910 when (BITSEL_u8_u1_1646_wire(0) /=  '0') else IMA88_900;
    -- logger for split-operator MUX_1657_inst flow-through 
    process(IMB45_1658) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1657_inst:flowthrough inputs: " & " BITSEL_u8_u1_1654_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1654_wire) & " IMA91_930 = "& Convert_SLV_To_Hex_String(IMA91_930) & " IMA90_920 = "& Convert_SLV_To_Hex_String(IMA90_920) & " outputs:" & " IMB45_1658= "  & Convert_SLV_To_Hex_String(IMB45_1658));
      --
    end process; 
    -- flow-through select operator MUX_1657_inst
    IMB45_1658 <= IMA91_930 when (BITSEL_u8_u1_1654_wire(0) /=  '0') else IMA90_920;
    -- logger for split-operator MUX_1665_inst flow-through 
    process(IMB46_1666) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1665_inst:flowthrough inputs: " & " BITSEL_u8_u1_1662_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1662_wire) & " IMA93_950 = "& Convert_SLV_To_Hex_String(IMA93_950) & " IMA92_940 = "& Convert_SLV_To_Hex_String(IMA92_940) & " outputs:" & " IMB46_1666= "  & Convert_SLV_To_Hex_String(IMB46_1666));
      --
    end process; 
    -- flow-through select operator MUX_1665_inst
    IMB46_1666 <= IMA93_950 when (BITSEL_u8_u1_1662_wire(0) /=  '0') else IMA92_940;
    -- logger for split-operator MUX_1673_inst flow-through 
    process(IMB47_1674) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1673_inst:flowthrough inputs: " & " BITSEL_u8_u1_1670_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1670_wire) & " IMA95_970 = "& Convert_SLV_To_Hex_String(IMA95_970) & " IMA94_960 = "& Convert_SLV_To_Hex_String(IMA94_960) & " outputs:" & " IMB47_1674= "  & Convert_SLV_To_Hex_String(IMB47_1674));
      --
    end process; 
    -- flow-through select operator MUX_1673_inst
    IMB47_1674 <= IMA95_970 when (BITSEL_u8_u1_1670_wire(0) /=  '0') else IMA94_960;
    -- logger for split-operator MUX_1681_inst flow-through 
    process(IMB48_1682) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1681_inst:flowthrough inputs: " & " BITSEL_u8_u1_1678_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1678_wire) & " IMA97_990 = "& Convert_SLV_To_Hex_String(IMA97_990) & " IMA96_980 = "& Convert_SLV_To_Hex_String(IMA96_980) & " outputs:" & " IMB48_1682= "  & Convert_SLV_To_Hex_String(IMB48_1682));
      --
    end process; 
    -- flow-through select operator MUX_1681_inst
    IMB48_1682 <= IMA97_990 when (BITSEL_u8_u1_1678_wire(0) /=  '0') else IMA96_980;
    -- logger for split-operator MUX_1689_inst flow-through 
    process(IMB49_1690) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1689_inst:flowthrough inputs: " & " BITSEL_u8_u1_1686_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1686_wire) & " IMA99_1010 = "& Convert_SLV_To_Hex_String(IMA99_1010) & " IMA98_1000 = "& Convert_SLV_To_Hex_String(IMA98_1000) & " outputs:" & " IMB49_1690= "  & Convert_SLV_To_Hex_String(IMB49_1690));
      --
    end process; 
    -- flow-through select operator MUX_1689_inst
    IMB49_1690 <= IMA99_1010 when (BITSEL_u8_u1_1686_wire(0) /=  '0') else IMA98_1000;
    -- logger for split-operator MUX_1697_inst flow-through 
    process(IMB50_1698) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1697_inst:flowthrough inputs: " & " BITSEL_u8_u1_1694_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1694_wire) & " IMA101_1030 = "& Convert_SLV_To_Hex_String(IMA101_1030) & " IMA100_1020 = "& Convert_SLV_To_Hex_String(IMA100_1020) & " outputs:" & " IMB50_1698= "  & Convert_SLV_To_Hex_String(IMB50_1698));
      --
    end process; 
    -- flow-through select operator MUX_1697_inst
    IMB50_1698 <= IMA101_1030 when (BITSEL_u8_u1_1694_wire(0) /=  '0') else IMA100_1020;
    -- logger for split-operator MUX_169_inst flow-through 
    process(IMA15_170) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_169_inst:flowthrough inputs: " & " BITSEL_u8_u1_164_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_164_wire) & " type_cast_166_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_166_wire_constant) & " type_cast_168_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_168_wire_constant) & " outputs:" & " IMA15_170= "  & Convert_SLV_To_Hex_String(IMA15_170));
      --
    end process; 
    -- flow-through select operator MUX_169_inst
    IMA15_170 <= type_cast_166_wire_constant when (BITSEL_u8_u1_164_wire(0) /=  '0') else type_cast_168_wire_constant;
    -- logger for split-operator MUX_1705_inst flow-through 
    process(IMB51_1706) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1705_inst:flowthrough inputs: " & " BITSEL_u8_u1_1702_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1702_wire) & " IMA103_1050 = "& Convert_SLV_To_Hex_String(IMA103_1050) & " IMA102_1040 = "& Convert_SLV_To_Hex_String(IMA102_1040) & " outputs:" & " IMB51_1706= "  & Convert_SLV_To_Hex_String(IMB51_1706));
      --
    end process; 
    -- flow-through select operator MUX_1705_inst
    IMB51_1706 <= IMA103_1050 when (BITSEL_u8_u1_1702_wire(0) /=  '0') else IMA102_1040;
    -- logger for split-operator MUX_1713_inst flow-through 
    process(IMB52_1714) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1713_inst:flowthrough inputs: " & " BITSEL_u8_u1_1710_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1710_wire) & " IMA105_1070 = "& Convert_SLV_To_Hex_String(IMA105_1070) & " IMA104_1060 = "& Convert_SLV_To_Hex_String(IMA104_1060) & " outputs:" & " IMB52_1714= "  & Convert_SLV_To_Hex_String(IMB52_1714));
      --
    end process; 
    -- flow-through select operator MUX_1713_inst
    IMB52_1714 <= IMA105_1070 when (BITSEL_u8_u1_1710_wire(0) /=  '0') else IMA104_1060;
    -- logger for split-operator MUX_1721_inst flow-through 
    process(IMB53_1722) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1721_inst:flowthrough inputs: " & " BITSEL_u8_u1_1718_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1718_wire) & " IMA107_1090 = "& Convert_SLV_To_Hex_String(IMA107_1090) & " IMA106_1080 = "& Convert_SLV_To_Hex_String(IMA106_1080) & " outputs:" & " IMB53_1722= "  & Convert_SLV_To_Hex_String(IMB53_1722));
      --
    end process; 
    -- flow-through select operator MUX_1721_inst
    IMB53_1722 <= IMA107_1090 when (BITSEL_u8_u1_1718_wire(0) /=  '0') else IMA106_1080;
    -- logger for split-operator MUX_1729_inst flow-through 
    process(IMB54_1730) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1729_inst:flowthrough inputs: " & " BITSEL_u8_u1_1726_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1726_wire) & " IMA109_1110 = "& Convert_SLV_To_Hex_String(IMA109_1110) & " IMA108_1100 = "& Convert_SLV_To_Hex_String(IMA108_1100) & " outputs:" & " IMB54_1730= "  & Convert_SLV_To_Hex_String(IMB54_1730));
      --
    end process; 
    -- flow-through select operator MUX_1729_inst
    IMB54_1730 <= IMA109_1110 when (BITSEL_u8_u1_1726_wire(0) /=  '0') else IMA108_1100;
    -- logger for split-operator MUX_1737_inst flow-through 
    process(IMB55_1738) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1737_inst:flowthrough inputs: " & " BITSEL_u8_u1_1734_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1734_wire) & " IMA111_1130 = "& Convert_SLV_To_Hex_String(IMA111_1130) & " IMA110_1120 = "& Convert_SLV_To_Hex_String(IMA110_1120) & " outputs:" & " IMB55_1738= "  & Convert_SLV_To_Hex_String(IMB55_1738));
      --
    end process; 
    -- flow-through select operator MUX_1737_inst
    IMB55_1738 <= IMA111_1130 when (BITSEL_u8_u1_1734_wire(0) /=  '0') else IMA110_1120;
    -- logger for split-operator MUX_1745_inst flow-through 
    process(IMB56_1746) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1745_inst:flowthrough inputs: " & " BITSEL_u8_u1_1742_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1742_wire) & " IMA113_1150 = "& Convert_SLV_To_Hex_String(IMA113_1150) & " IMA112_1140 = "& Convert_SLV_To_Hex_String(IMA112_1140) & " outputs:" & " IMB56_1746= "  & Convert_SLV_To_Hex_String(IMB56_1746));
      --
    end process; 
    -- flow-through select operator MUX_1745_inst
    IMB56_1746 <= IMA113_1150 when (BITSEL_u8_u1_1742_wire(0) /=  '0') else IMA112_1140;
    -- logger for split-operator MUX_1753_inst flow-through 
    process(IMB57_1754) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1753_inst:flowthrough inputs: " & " BITSEL_u8_u1_1750_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1750_wire) & " IMA115_1170 = "& Convert_SLV_To_Hex_String(IMA115_1170) & " IMA114_1160 = "& Convert_SLV_To_Hex_String(IMA114_1160) & " outputs:" & " IMB57_1754= "  & Convert_SLV_To_Hex_String(IMB57_1754));
      --
    end process; 
    -- flow-through select operator MUX_1753_inst
    IMB57_1754 <= IMA115_1170 when (BITSEL_u8_u1_1750_wire(0) /=  '0') else IMA114_1160;
    -- logger for split-operator MUX_1761_inst flow-through 
    process(IMB58_1762) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1761_inst:flowthrough inputs: " & " BITSEL_u8_u1_1758_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1758_wire) & " IMA117_1190 = "& Convert_SLV_To_Hex_String(IMA117_1190) & " IMA116_1180 = "& Convert_SLV_To_Hex_String(IMA116_1180) & " outputs:" & " IMB58_1762= "  & Convert_SLV_To_Hex_String(IMB58_1762));
      --
    end process; 
    -- flow-through select operator MUX_1761_inst
    IMB58_1762 <= IMA117_1190 when (BITSEL_u8_u1_1758_wire(0) /=  '0') else IMA116_1180;
    -- logger for split-operator MUX_1769_inst flow-through 
    process(IMB59_1770) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1769_inst:flowthrough inputs: " & " BITSEL_u8_u1_1766_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1766_wire) & " IMA119_1210 = "& Convert_SLV_To_Hex_String(IMA119_1210) & " IMA118_1200 = "& Convert_SLV_To_Hex_String(IMA118_1200) & " outputs:" & " IMB59_1770= "  & Convert_SLV_To_Hex_String(IMB59_1770));
      --
    end process; 
    -- flow-through select operator MUX_1769_inst
    IMB59_1770 <= IMA119_1210 when (BITSEL_u8_u1_1766_wire(0) /=  '0') else IMA118_1200;
    -- logger for split-operator MUX_1777_inst flow-through 
    process(IMB60_1778) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1777_inst:flowthrough inputs: " & " BITSEL_u8_u1_1774_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1774_wire) & " IMA121_1230 = "& Convert_SLV_To_Hex_String(IMA121_1230) & " IMA120_1220 = "& Convert_SLV_To_Hex_String(IMA120_1220) & " outputs:" & " IMB60_1778= "  & Convert_SLV_To_Hex_String(IMB60_1778));
      --
    end process; 
    -- flow-through select operator MUX_1777_inst
    IMB60_1778 <= IMA121_1230 when (BITSEL_u8_u1_1774_wire(0) /=  '0') else IMA120_1220;
    -- logger for split-operator MUX_1785_inst flow-through 
    process(IMB61_1786) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1785_inst:flowthrough inputs: " & " BITSEL_u8_u1_1782_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1782_wire) & " IMA123_1250 = "& Convert_SLV_To_Hex_String(IMA123_1250) & " IMA122_1240 = "& Convert_SLV_To_Hex_String(IMA122_1240) & " outputs:" & " IMB61_1786= "  & Convert_SLV_To_Hex_String(IMB61_1786));
      --
    end process; 
    -- flow-through select operator MUX_1785_inst
    IMB61_1786 <= IMA123_1250 when (BITSEL_u8_u1_1782_wire(0) /=  '0') else IMA122_1240;
    -- logger for split-operator MUX_1793_inst flow-through 
    process(IMB62_1794) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1793_inst:flowthrough inputs: " & " BITSEL_u8_u1_1790_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1790_wire) & " IMA125_1270 = "& Convert_SLV_To_Hex_String(IMA125_1270) & " IMA124_1260 = "& Convert_SLV_To_Hex_String(IMA124_1260) & " outputs:" & " IMB62_1794= "  & Convert_SLV_To_Hex_String(IMB62_1794));
      --
    end process; 
    -- flow-through select operator MUX_1793_inst
    IMB62_1794 <= IMA125_1270 when (BITSEL_u8_u1_1790_wire(0) /=  '0') else IMA124_1260;
    -- logger for split-operator MUX_179_inst flow-through 
    process(IMA16_180) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_179_inst:flowthrough inputs: " & " BITSEL_u8_u1_174_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_174_wire) & " type_cast_176_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_176_wire_constant) & " type_cast_178_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_178_wire_constant) & " outputs:" & " IMA16_180= "  & Convert_SLV_To_Hex_String(IMA16_180));
      --
    end process; 
    -- flow-through select operator MUX_179_inst
    IMA16_180 <= type_cast_176_wire_constant when (BITSEL_u8_u1_174_wire(0) /=  '0') else type_cast_178_wire_constant;
    -- logger for split-operator MUX_1801_inst flow-through 
    process(IMB63_1802) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1801_inst:flowthrough inputs: " & " BITSEL_u8_u1_1798_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1798_wire) & " IMA127_1290 = "& Convert_SLV_To_Hex_String(IMA127_1290) & " IMA126_1280 = "& Convert_SLV_To_Hex_String(IMA126_1280) & " outputs:" & " IMB63_1802= "  & Convert_SLV_To_Hex_String(IMB63_1802));
      --
    end process; 
    -- flow-through select operator MUX_1801_inst
    IMB63_1802 <= IMA127_1290 when (BITSEL_u8_u1_1798_wire(0) /=  '0') else IMA126_1280;
    -- logger for split-operator MUX_1809_inst flow-through 
    process(IMC0_1810) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1809_inst:flowthrough inputs: " & " BITSEL_u8_u1_1806_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1806_wire) & " IMB1_1306 = "& Convert_SLV_To_Hex_String(IMB1_1306) & " IMB0_1298 = "& Convert_SLV_To_Hex_String(IMB0_1298) & " outputs:" & " IMC0_1810= "  & Convert_SLV_To_Hex_String(IMC0_1810));
      --
    end process; 
    -- flow-through select operator MUX_1809_inst
    IMC0_1810 <= IMB1_1306 when (BITSEL_u8_u1_1806_wire(0) /=  '0') else IMB0_1298;
    -- logger for split-operator MUX_1817_inst flow-through 
    process(IMC1_1818) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1817_inst:flowthrough inputs: " & " BITSEL_u8_u1_1814_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1814_wire) & " IMB3_1322 = "& Convert_SLV_To_Hex_String(IMB3_1322) & " IMB2_1314 = "& Convert_SLV_To_Hex_String(IMB2_1314) & " outputs:" & " IMC1_1818= "  & Convert_SLV_To_Hex_String(IMC1_1818));
      --
    end process; 
    -- flow-through select operator MUX_1817_inst
    IMC1_1818 <= IMB3_1322 when (BITSEL_u8_u1_1814_wire(0) /=  '0') else IMB2_1314;
    -- logger for split-operator MUX_1825_inst flow-through 
    process(IMC2_1826) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1825_inst:flowthrough inputs: " & " BITSEL_u8_u1_1822_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1822_wire) & " IMB5_1338 = "& Convert_SLV_To_Hex_String(IMB5_1338) & " IMB4_1330 = "& Convert_SLV_To_Hex_String(IMB4_1330) & " outputs:" & " IMC2_1826= "  & Convert_SLV_To_Hex_String(IMC2_1826));
      --
    end process; 
    -- flow-through select operator MUX_1825_inst
    IMC2_1826 <= IMB5_1338 when (BITSEL_u8_u1_1822_wire(0) /=  '0') else IMB4_1330;
    -- logger for split-operator MUX_1833_inst flow-through 
    process(IMC3_1834) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1833_inst:flowthrough inputs: " & " BITSEL_u8_u1_1830_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1830_wire) & " IMB7_1354 = "& Convert_SLV_To_Hex_String(IMB7_1354) & " IMB6_1346 = "& Convert_SLV_To_Hex_String(IMB6_1346) & " outputs:" & " IMC3_1834= "  & Convert_SLV_To_Hex_String(IMC3_1834));
      --
    end process; 
    -- flow-through select operator MUX_1833_inst
    IMC3_1834 <= IMB7_1354 when (BITSEL_u8_u1_1830_wire(0) /=  '0') else IMB6_1346;
    -- logger for split-operator MUX_1841_inst flow-through 
    process(IMC4_1842) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1841_inst:flowthrough inputs: " & " BITSEL_u8_u1_1838_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1838_wire) & " IMB9_1370 = "& Convert_SLV_To_Hex_String(IMB9_1370) & " IMB8_1362 = "& Convert_SLV_To_Hex_String(IMB8_1362) & " outputs:" & " IMC4_1842= "  & Convert_SLV_To_Hex_String(IMC4_1842));
      --
    end process; 
    -- flow-through select operator MUX_1841_inst
    IMC4_1842 <= IMB9_1370 when (BITSEL_u8_u1_1838_wire(0) /=  '0') else IMB8_1362;
    -- logger for split-operator MUX_1849_inst flow-through 
    process(IMC5_1850) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1849_inst:flowthrough inputs: " & " BITSEL_u8_u1_1846_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1846_wire) & " IMB11_1386 = "& Convert_SLV_To_Hex_String(IMB11_1386) & " IMB10_1378 = "& Convert_SLV_To_Hex_String(IMB10_1378) & " outputs:" & " IMC5_1850= "  & Convert_SLV_To_Hex_String(IMC5_1850));
      --
    end process; 
    -- flow-through select operator MUX_1849_inst
    IMC5_1850 <= IMB11_1386 when (BITSEL_u8_u1_1846_wire(0) /=  '0') else IMB10_1378;
    -- logger for split-operator MUX_1857_inst flow-through 
    process(IMC6_1858) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1857_inst:flowthrough inputs: " & " BITSEL_u8_u1_1854_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1854_wire) & " IMB13_1402 = "& Convert_SLV_To_Hex_String(IMB13_1402) & " IMB12_1394 = "& Convert_SLV_To_Hex_String(IMB12_1394) & " outputs:" & " IMC6_1858= "  & Convert_SLV_To_Hex_String(IMC6_1858));
      --
    end process; 
    -- flow-through select operator MUX_1857_inst
    IMC6_1858 <= IMB13_1402 when (BITSEL_u8_u1_1854_wire(0) /=  '0') else IMB12_1394;
    -- logger for split-operator MUX_1865_inst flow-through 
    process(IMC7_1866) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1865_inst:flowthrough inputs: " & " BITSEL_u8_u1_1862_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1862_wire) & " IMB15_1418 = "& Convert_SLV_To_Hex_String(IMB15_1418) & " IMB14_1410 = "& Convert_SLV_To_Hex_String(IMB14_1410) & " outputs:" & " IMC7_1866= "  & Convert_SLV_To_Hex_String(IMC7_1866));
      --
    end process; 
    -- flow-through select operator MUX_1865_inst
    IMC7_1866 <= IMB15_1418 when (BITSEL_u8_u1_1862_wire(0) /=  '0') else IMB14_1410;
    -- logger for split-operator MUX_1873_inst flow-through 
    process(IMC8_1874) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1873_inst:flowthrough inputs: " & " BITSEL_u8_u1_1870_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1870_wire) & " IMB17_1434 = "& Convert_SLV_To_Hex_String(IMB17_1434) & " IMB16_1426 = "& Convert_SLV_To_Hex_String(IMB16_1426) & " outputs:" & " IMC8_1874= "  & Convert_SLV_To_Hex_String(IMC8_1874));
      --
    end process; 
    -- flow-through select operator MUX_1873_inst
    IMC8_1874 <= IMB17_1434 when (BITSEL_u8_u1_1870_wire(0) /=  '0') else IMB16_1426;
    -- logger for split-operator MUX_1881_inst flow-through 
    process(IMC9_1882) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1881_inst:flowthrough inputs: " & " BITSEL_u8_u1_1878_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1878_wire) & " IMB19_1450 = "& Convert_SLV_To_Hex_String(IMB19_1450) & " IMB18_1442 = "& Convert_SLV_To_Hex_String(IMB18_1442) & " outputs:" & " IMC9_1882= "  & Convert_SLV_To_Hex_String(IMC9_1882));
      --
    end process; 
    -- flow-through select operator MUX_1881_inst
    IMC9_1882 <= IMB19_1450 when (BITSEL_u8_u1_1878_wire(0) /=  '0') else IMB18_1442;
    -- logger for split-operator MUX_1889_inst flow-through 
    process(IMC10_1890) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1889_inst:flowthrough inputs: " & " BITSEL_u8_u1_1886_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1886_wire) & " IMB21_1466 = "& Convert_SLV_To_Hex_String(IMB21_1466) & " IMB20_1458 = "& Convert_SLV_To_Hex_String(IMB20_1458) & " outputs:" & " IMC10_1890= "  & Convert_SLV_To_Hex_String(IMC10_1890));
      --
    end process; 
    -- flow-through select operator MUX_1889_inst
    IMC10_1890 <= IMB21_1466 when (BITSEL_u8_u1_1886_wire(0) /=  '0') else IMB20_1458;
    -- logger for split-operator MUX_1897_inst flow-through 
    process(IMC11_1898) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1897_inst:flowthrough inputs: " & " BITSEL_u8_u1_1894_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1894_wire) & " IMB23_1482 = "& Convert_SLV_To_Hex_String(IMB23_1482) & " IMB22_1474 = "& Convert_SLV_To_Hex_String(IMB22_1474) & " outputs:" & " IMC11_1898= "  & Convert_SLV_To_Hex_String(IMC11_1898));
      --
    end process; 
    -- flow-through select operator MUX_1897_inst
    IMC11_1898 <= IMB23_1482 when (BITSEL_u8_u1_1894_wire(0) /=  '0') else IMB22_1474;
    -- logger for split-operator MUX_189_inst flow-through 
    process(IMA17_190) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_189_inst:flowthrough inputs: " & " BITSEL_u8_u1_184_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_184_wire) & " type_cast_186_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_186_wire_constant) & " type_cast_188_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_188_wire_constant) & " outputs:" & " IMA17_190= "  & Convert_SLV_To_Hex_String(IMA17_190));
      --
    end process; 
    -- flow-through select operator MUX_189_inst
    IMA17_190 <= type_cast_186_wire_constant when (BITSEL_u8_u1_184_wire(0) /=  '0') else type_cast_188_wire_constant;
    -- logger for split-operator MUX_1905_inst flow-through 
    process(IMC12_1906) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1905_inst:flowthrough inputs: " & " BITSEL_u8_u1_1902_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1902_wire) & " IMB25_1498 = "& Convert_SLV_To_Hex_String(IMB25_1498) & " IMB24_1490 = "& Convert_SLV_To_Hex_String(IMB24_1490) & " outputs:" & " IMC12_1906= "  & Convert_SLV_To_Hex_String(IMC12_1906));
      --
    end process; 
    -- flow-through select operator MUX_1905_inst
    IMC12_1906 <= IMB25_1498 when (BITSEL_u8_u1_1902_wire(0) /=  '0') else IMB24_1490;
    -- logger for split-operator MUX_1913_inst flow-through 
    process(IMC13_1914) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1913_inst:flowthrough inputs: " & " BITSEL_u8_u1_1910_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1910_wire) & " IMB27_1514 = "& Convert_SLV_To_Hex_String(IMB27_1514) & " IMB26_1506 = "& Convert_SLV_To_Hex_String(IMB26_1506) & " outputs:" & " IMC13_1914= "  & Convert_SLV_To_Hex_String(IMC13_1914));
      --
    end process; 
    -- flow-through select operator MUX_1913_inst
    IMC13_1914 <= IMB27_1514 when (BITSEL_u8_u1_1910_wire(0) /=  '0') else IMB26_1506;
    -- logger for split-operator MUX_1921_inst flow-through 
    process(IMC14_1922) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1921_inst:flowthrough inputs: " & " BITSEL_u8_u1_1918_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1918_wire) & " IMB29_1530 = "& Convert_SLV_To_Hex_String(IMB29_1530) & " IMB28_1522 = "& Convert_SLV_To_Hex_String(IMB28_1522) & " outputs:" & " IMC14_1922= "  & Convert_SLV_To_Hex_String(IMC14_1922));
      --
    end process; 
    -- flow-through select operator MUX_1921_inst
    IMC14_1922 <= IMB29_1530 when (BITSEL_u8_u1_1918_wire(0) /=  '0') else IMB28_1522;
    -- logger for split-operator MUX_1929_inst flow-through 
    process(IMC15_1930) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1929_inst:flowthrough inputs: " & " BITSEL_u8_u1_1926_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1926_wire) & " IMB31_1546 = "& Convert_SLV_To_Hex_String(IMB31_1546) & " IMB30_1538 = "& Convert_SLV_To_Hex_String(IMB30_1538) & " outputs:" & " IMC15_1930= "  & Convert_SLV_To_Hex_String(IMC15_1930));
      --
    end process; 
    -- flow-through select operator MUX_1929_inst
    IMC15_1930 <= IMB31_1546 when (BITSEL_u8_u1_1926_wire(0) /=  '0') else IMB30_1538;
    -- logger for split-operator MUX_1937_inst flow-through 
    process(IMC16_1938) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1937_inst:flowthrough inputs: " & " BITSEL_u8_u1_1934_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1934_wire) & " IMB33_1562 = "& Convert_SLV_To_Hex_String(IMB33_1562) & " IMB32_1554 = "& Convert_SLV_To_Hex_String(IMB32_1554) & " outputs:" & " IMC16_1938= "  & Convert_SLV_To_Hex_String(IMC16_1938));
      --
    end process; 
    -- flow-through select operator MUX_1937_inst
    IMC16_1938 <= IMB33_1562 when (BITSEL_u8_u1_1934_wire(0) /=  '0') else IMB32_1554;
    -- logger for split-operator MUX_1945_inst flow-through 
    process(IMC17_1946) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1945_inst:flowthrough inputs: " & " BITSEL_u8_u1_1942_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1942_wire) & " IMB35_1578 = "& Convert_SLV_To_Hex_String(IMB35_1578) & " IMB34_1570 = "& Convert_SLV_To_Hex_String(IMB34_1570) & " outputs:" & " IMC17_1946= "  & Convert_SLV_To_Hex_String(IMC17_1946));
      --
    end process; 
    -- flow-through select operator MUX_1945_inst
    IMC17_1946 <= IMB35_1578 when (BITSEL_u8_u1_1942_wire(0) /=  '0') else IMB34_1570;
    -- logger for split-operator MUX_1953_inst flow-through 
    process(IMC18_1954) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1953_inst:flowthrough inputs: " & " BITSEL_u8_u1_1950_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1950_wire) & " IMB37_1594 = "& Convert_SLV_To_Hex_String(IMB37_1594) & " IMB36_1586 = "& Convert_SLV_To_Hex_String(IMB36_1586) & " outputs:" & " IMC18_1954= "  & Convert_SLV_To_Hex_String(IMC18_1954));
      --
    end process; 
    -- flow-through select operator MUX_1953_inst
    IMC18_1954 <= IMB37_1594 when (BITSEL_u8_u1_1950_wire(0) /=  '0') else IMB36_1586;
    -- logger for split-operator MUX_1961_inst flow-through 
    process(IMC19_1962) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1961_inst:flowthrough inputs: " & " BITSEL_u8_u1_1958_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1958_wire) & " IMB39_1610 = "& Convert_SLV_To_Hex_String(IMB39_1610) & " IMB38_1602 = "& Convert_SLV_To_Hex_String(IMB38_1602) & " outputs:" & " IMC19_1962= "  & Convert_SLV_To_Hex_String(IMC19_1962));
      --
    end process; 
    -- flow-through select operator MUX_1961_inst
    IMC19_1962 <= IMB39_1610 when (BITSEL_u8_u1_1958_wire(0) /=  '0') else IMB38_1602;
    -- logger for split-operator MUX_1969_inst flow-through 
    process(IMC20_1970) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1969_inst:flowthrough inputs: " & " BITSEL_u8_u1_1966_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1966_wire) & " IMB41_1626 = "& Convert_SLV_To_Hex_String(IMB41_1626) & " IMB40_1618 = "& Convert_SLV_To_Hex_String(IMB40_1618) & " outputs:" & " IMC20_1970= "  & Convert_SLV_To_Hex_String(IMC20_1970));
      --
    end process; 
    -- flow-through select operator MUX_1969_inst
    IMC20_1970 <= IMB41_1626 when (BITSEL_u8_u1_1966_wire(0) /=  '0') else IMB40_1618;
    -- logger for split-operator MUX_1977_inst flow-through 
    process(IMC21_1978) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1977_inst:flowthrough inputs: " & " BITSEL_u8_u1_1974_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1974_wire) & " IMB43_1642 = "& Convert_SLV_To_Hex_String(IMB43_1642) & " IMB42_1634 = "& Convert_SLV_To_Hex_String(IMB42_1634) & " outputs:" & " IMC21_1978= "  & Convert_SLV_To_Hex_String(IMC21_1978));
      --
    end process; 
    -- flow-through select operator MUX_1977_inst
    IMC21_1978 <= IMB43_1642 when (BITSEL_u8_u1_1974_wire(0) /=  '0') else IMB42_1634;
    -- logger for split-operator MUX_1985_inst flow-through 
    process(IMC22_1986) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1985_inst:flowthrough inputs: " & " BITSEL_u8_u1_1982_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1982_wire) & " IMB45_1658 = "& Convert_SLV_To_Hex_String(IMB45_1658) & " IMB44_1650 = "& Convert_SLV_To_Hex_String(IMB44_1650) & " outputs:" & " IMC22_1986= "  & Convert_SLV_To_Hex_String(IMC22_1986));
      --
    end process; 
    -- flow-through select operator MUX_1985_inst
    IMC22_1986 <= IMB45_1658 when (BITSEL_u8_u1_1982_wire(0) /=  '0') else IMB44_1650;
    -- logger for split-operator MUX_1993_inst flow-through 
    process(IMC23_1994) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_1993_inst:flowthrough inputs: " & " BITSEL_u8_u1_1990_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1990_wire) & " IMB47_1674 = "& Convert_SLV_To_Hex_String(IMB47_1674) & " IMB46_1666 = "& Convert_SLV_To_Hex_String(IMB46_1666) & " outputs:" & " IMC23_1994= "  & Convert_SLV_To_Hex_String(IMC23_1994));
      --
    end process; 
    -- flow-through select operator MUX_1993_inst
    IMC23_1994 <= IMB47_1674 when (BITSEL_u8_u1_1990_wire(0) /=  '0') else IMB46_1666;
    -- logger for split-operator MUX_199_inst flow-through 
    process(IMA18_200) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_199_inst:flowthrough inputs: " & " BITSEL_u8_u1_194_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_194_wire) & " type_cast_196_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_196_wire_constant) & " type_cast_198_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_198_wire_constant) & " outputs:" & " IMA18_200= "  & Convert_SLV_To_Hex_String(IMA18_200));
      --
    end process; 
    -- flow-through select operator MUX_199_inst
    IMA18_200 <= type_cast_196_wire_constant when (BITSEL_u8_u1_194_wire(0) /=  '0') else type_cast_198_wire_constant;
    -- logger for split-operator MUX_19_inst flow-through 
    process(IMA0_20) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_19_inst:flowthrough inputs: " & " BITSEL_u8_u1_13_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_13_wire) & " type_cast_16_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_16_wire_constant) & " type_cast_18_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_18_wire_constant) & " outputs:" & " IMA0_20= "  & Convert_SLV_To_Hex_String(IMA0_20));
      --
    end process; 
    -- flow-through select operator MUX_19_inst
    IMA0_20 <= type_cast_16_wire_constant when (BITSEL_u8_u1_13_wire(0) /=  '0') else type_cast_18_wire_constant;
    -- logger for split-operator MUX_2001_inst flow-through 
    process(IMC24_2002) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_2001_inst:flowthrough inputs: " & " BITSEL_u8_u1_1998_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1998_wire) & " IMB49_1690 = "& Convert_SLV_To_Hex_String(IMB49_1690) & " IMB48_1682 = "& Convert_SLV_To_Hex_String(IMB48_1682) & " outputs:" & " IMC24_2002= "  & Convert_SLV_To_Hex_String(IMC24_2002));
      --
    end process; 
    -- flow-through select operator MUX_2001_inst
    IMC24_2002 <= IMB49_1690 when (BITSEL_u8_u1_1998_wire(0) /=  '0') else IMB48_1682;
    -- logger for split-operator MUX_2009_inst flow-through 
    process(IMC25_2010) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_2009_inst:flowthrough inputs: " & " BITSEL_u8_u1_2006_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_2006_wire) & " IMB51_1706 = "& Convert_SLV_To_Hex_String(IMB51_1706) & " IMB50_1698 = "& Convert_SLV_To_Hex_String(IMB50_1698) & " outputs:" & " IMC25_2010= "  & Convert_SLV_To_Hex_String(IMC25_2010));
      --
    end process; 
    -- flow-through select operator MUX_2009_inst
    IMC25_2010 <= IMB51_1706 when (BITSEL_u8_u1_2006_wire(0) /=  '0') else IMB50_1698;
    -- logger for split-operator MUX_2017_inst flow-through 
    process(IMC26_2018) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_2017_inst:flowthrough inputs: " & " BITSEL_u8_u1_2014_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_2014_wire) & " IMB53_1722 = "& Convert_SLV_To_Hex_String(IMB53_1722) & " IMB52_1714 = "& Convert_SLV_To_Hex_String(IMB52_1714) & " outputs:" & " IMC26_2018= "  & Convert_SLV_To_Hex_String(IMC26_2018));
      --
    end process; 
    -- flow-through select operator MUX_2017_inst
    IMC26_2018 <= IMB53_1722 when (BITSEL_u8_u1_2014_wire(0) /=  '0') else IMB52_1714;
    -- logger for split-operator MUX_2025_inst flow-through 
    process(IMC27_2026) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_2025_inst:flowthrough inputs: " & " BITSEL_u8_u1_2022_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_2022_wire) & " IMB55_1738 = "& Convert_SLV_To_Hex_String(IMB55_1738) & " IMB54_1730 = "& Convert_SLV_To_Hex_String(IMB54_1730) & " outputs:" & " IMC27_2026= "  & Convert_SLV_To_Hex_String(IMC27_2026));
      --
    end process; 
    -- flow-through select operator MUX_2025_inst
    IMC27_2026 <= IMB55_1738 when (BITSEL_u8_u1_2022_wire(0) /=  '0') else IMB54_1730;
    -- logger for split-operator MUX_2033_inst flow-through 
    process(IMC28_2034) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_2033_inst:flowthrough inputs: " & " BITSEL_u8_u1_2030_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_2030_wire) & " IMB57_1754 = "& Convert_SLV_To_Hex_String(IMB57_1754) & " IMB56_1746 = "& Convert_SLV_To_Hex_String(IMB56_1746) & " outputs:" & " IMC28_2034= "  & Convert_SLV_To_Hex_String(IMC28_2034));
      --
    end process; 
    -- flow-through select operator MUX_2033_inst
    IMC28_2034 <= IMB57_1754 when (BITSEL_u8_u1_2030_wire(0) /=  '0') else IMB56_1746;
    -- logger for split-operator MUX_2041_inst flow-through 
    process(IMC29_2042) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_2041_inst:flowthrough inputs: " & " BITSEL_u8_u1_2038_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_2038_wire) & " IMB59_1770 = "& Convert_SLV_To_Hex_String(IMB59_1770) & " IMB58_1762 = "& Convert_SLV_To_Hex_String(IMB58_1762) & " outputs:" & " IMC29_2042= "  & Convert_SLV_To_Hex_String(IMC29_2042));
      --
    end process; 
    -- flow-through select operator MUX_2041_inst
    IMC29_2042 <= IMB59_1770 when (BITSEL_u8_u1_2038_wire(0) /=  '0') else IMB58_1762;
    -- logger for split-operator MUX_2049_inst flow-through 
    process(IMC30_2050) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_2049_inst:flowthrough inputs: " & " BITSEL_u8_u1_2046_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_2046_wire) & " IMB61_1786 = "& Convert_SLV_To_Hex_String(IMB61_1786) & " IMB60_1778 = "& Convert_SLV_To_Hex_String(IMB60_1778) & " outputs:" & " IMC30_2050= "  & Convert_SLV_To_Hex_String(IMC30_2050));
      --
    end process; 
    -- flow-through select operator MUX_2049_inst
    IMC30_2050 <= IMB61_1786 when (BITSEL_u8_u1_2046_wire(0) /=  '0') else IMB60_1778;
    -- logger for split-operator MUX_2057_inst flow-through 
    process(IMC31_2058) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_2057_inst:flowthrough inputs: " & " BITSEL_u8_u1_2054_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_2054_wire) & " IMB63_1802 = "& Convert_SLV_To_Hex_String(IMB63_1802) & " IMB62_1794 = "& Convert_SLV_To_Hex_String(IMB62_1794) & " outputs:" & " IMC31_2058= "  & Convert_SLV_To_Hex_String(IMC31_2058));
      --
    end process; 
    -- flow-through select operator MUX_2057_inst
    IMC31_2058 <= IMB63_1802 when (BITSEL_u8_u1_2054_wire(0) /=  '0') else IMB62_1794;
    -- logger for split-operator MUX_2065_inst flow-through 
    process(IMD0_2066) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_2065_inst:flowthrough inputs: " & " BITSEL_u8_u1_2062_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_2062_wire) & " IMC1_1818 = "& Convert_SLV_To_Hex_String(IMC1_1818) & " IMC0_1810 = "& Convert_SLV_To_Hex_String(IMC0_1810) & " outputs:" & " IMD0_2066= "  & Convert_SLV_To_Hex_String(IMD0_2066));
      --
    end process; 
    -- flow-through select operator MUX_2065_inst
    IMD0_2066 <= IMC1_1818 when (BITSEL_u8_u1_2062_wire(0) /=  '0') else IMC0_1810;
    -- logger for split-operator MUX_2073_inst flow-through 
    process(IMD1_2074) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_2073_inst:flowthrough inputs: " & " BITSEL_u8_u1_2070_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_2070_wire) & " IMC3_1834 = "& Convert_SLV_To_Hex_String(IMC3_1834) & " IMC2_1826 = "& Convert_SLV_To_Hex_String(IMC2_1826) & " outputs:" & " IMD1_2074= "  & Convert_SLV_To_Hex_String(IMD1_2074));
      --
    end process; 
    -- flow-through select operator MUX_2073_inst
    IMD1_2074 <= IMC3_1834 when (BITSEL_u8_u1_2070_wire(0) /=  '0') else IMC2_1826;
    -- logger for split-operator MUX_2081_inst flow-through 
    process(IMD2_2082) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_2081_inst:flowthrough inputs: " & " BITSEL_u8_u1_2078_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_2078_wire) & " IMC5_1850 = "& Convert_SLV_To_Hex_String(IMC5_1850) & " IMC4_1842 = "& Convert_SLV_To_Hex_String(IMC4_1842) & " outputs:" & " IMD2_2082= "  & Convert_SLV_To_Hex_String(IMD2_2082));
      --
    end process; 
    -- flow-through select operator MUX_2081_inst
    IMD2_2082 <= IMC5_1850 when (BITSEL_u8_u1_2078_wire(0) /=  '0') else IMC4_1842;
    -- logger for split-operator MUX_2089_inst flow-through 
    process(IMD3_2090) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_2089_inst:flowthrough inputs: " & " BITSEL_u8_u1_2086_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_2086_wire) & " IMC7_1866 = "& Convert_SLV_To_Hex_String(IMC7_1866) & " IMC6_1858 = "& Convert_SLV_To_Hex_String(IMC6_1858) & " outputs:" & " IMD3_2090= "  & Convert_SLV_To_Hex_String(IMD3_2090));
      --
    end process; 
    -- flow-through select operator MUX_2089_inst
    IMD3_2090 <= IMC7_1866 when (BITSEL_u8_u1_2086_wire(0) /=  '0') else IMC6_1858;
    -- logger for split-operator MUX_2097_inst flow-through 
    process(IMD4_2098) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_2097_inst:flowthrough inputs: " & " BITSEL_u8_u1_2094_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_2094_wire) & " IMC9_1882 = "& Convert_SLV_To_Hex_String(IMC9_1882) & " IMC8_1874 = "& Convert_SLV_To_Hex_String(IMC8_1874) & " outputs:" & " IMD4_2098= "  & Convert_SLV_To_Hex_String(IMD4_2098));
      --
    end process; 
    -- flow-through select operator MUX_2097_inst
    IMD4_2098 <= IMC9_1882 when (BITSEL_u8_u1_2094_wire(0) /=  '0') else IMC8_1874;
    -- logger for split-operator MUX_209_inst flow-through 
    process(IMA19_210) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_209_inst:flowthrough inputs: " & " BITSEL_u8_u1_204_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_204_wire) & " type_cast_206_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_206_wire_constant) & " type_cast_208_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_208_wire_constant) & " outputs:" & " IMA19_210= "  & Convert_SLV_To_Hex_String(IMA19_210));
      --
    end process; 
    -- flow-through select operator MUX_209_inst
    IMA19_210 <= type_cast_206_wire_constant when (BITSEL_u8_u1_204_wire(0) /=  '0') else type_cast_208_wire_constant;
    -- logger for split-operator MUX_2105_inst flow-through 
    process(IMD5_2106) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_2105_inst:flowthrough inputs: " & " BITSEL_u8_u1_2102_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_2102_wire) & " IMC11_1898 = "& Convert_SLV_To_Hex_String(IMC11_1898) & " IMC10_1890 = "& Convert_SLV_To_Hex_String(IMC10_1890) & " outputs:" & " IMD5_2106= "  & Convert_SLV_To_Hex_String(IMD5_2106));
      --
    end process; 
    -- flow-through select operator MUX_2105_inst
    IMD5_2106 <= IMC11_1898 when (BITSEL_u8_u1_2102_wire(0) /=  '0') else IMC10_1890;
    -- logger for split-operator MUX_2113_inst flow-through 
    process(IMD6_2114) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_2113_inst:flowthrough inputs: " & " BITSEL_u8_u1_2110_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_2110_wire) & " IMC13_1914 = "& Convert_SLV_To_Hex_String(IMC13_1914) & " IMC12_1906 = "& Convert_SLV_To_Hex_String(IMC12_1906) & " outputs:" & " IMD6_2114= "  & Convert_SLV_To_Hex_String(IMD6_2114));
      --
    end process; 
    -- flow-through select operator MUX_2113_inst
    IMD6_2114 <= IMC13_1914 when (BITSEL_u8_u1_2110_wire(0) /=  '0') else IMC12_1906;
    -- logger for split-operator MUX_2121_inst flow-through 
    process(IMD7_2122) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_2121_inst:flowthrough inputs: " & " BITSEL_u8_u1_2118_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_2118_wire) & " IMC15_1930 = "& Convert_SLV_To_Hex_String(IMC15_1930) & " IMC14_1922 = "& Convert_SLV_To_Hex_String(IMC14_1922) & " outputs:" & " IMD7_2122= "  & Convert_SLV_To_Hex_String(IMD7_2122));
      --
    end process; 
    -- flow-through select operator MUX_2121_inst
    IMD7_2122 <= IMC15_1930 when (BITSEL_u8_u1_2118_wire(0) /=  '0') else IMC14_1922;
    -- logger for split-operator MUX_2129_inst flow-through 
    process(IMD8_2130) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_2129_inst:flowthrough inputs: " & " BITSEL_u8_u1_2126_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_2126_wire) & " IMC17_1946 = "& Convert_SLV_To_Hex_String(IMC17_1946) & " IMC16_1938 = "& Convert_SLV_To_Hex_String(IMC16_1938) & " outputs:" & " IMD8_2130= "  & Convert_SLV_To_Hex_String(IMD8_2130));
      --
    end process; 
    -- flow-through select operator MUX_2129_inst
    IMD8_2130 <= IMC17_1946 when (BITSEL_u8_u1_2126_wire(0) /=  '0') else IMC16_1938;
    -- logger for split-operator MUX_2137_inst flow-through 
    process(IMD9_2138) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_2137_inst:flowthrough inputs: " & " BITSEL_u8_u1_2134_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_2134_wire) & " IMC19_1962 = "& Convert_SLV_To_Hex_String(IMC19_1962) & " IMC18_1954 = "& Convert_SLV_To_Hex_String(IMC18_1954) & " outputs:" & " IMD9_2138= "  & Convert_SLV_To_Hex_String(IMD9_2138));
      --
    end process; 
    -- flow-through select operator MUX_2137_inst
    IMD9_2138 <= IMC19_1962 when (BITSEL_u8_u1_2134_wire(0) /=  '0') else IMC18_1954;
    -- logger for split-operator MUX_2145_inst flow-through 
    process(IMD10_2146) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_2145_inst:flowthrough inputs: " & " BITSEL_u8_u1_2142_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_2142_wire) & " IMC21_1978 = "& Convert_SLV_To_Hex_String(IMC21_1978) & " IMC20_1970 = "& Convert_SLV_To_Hex_String(IMC20_1970) & " outputs:" & " IMD10_2146= "  & Convert_SLV_To_Hex_String(IMD10_2146));
      --
    end process; 
    -- flow-through select operator MUX_2145_inst
    IMD10_2146 <= IMC21_1978 when (BITSEL_u8_u1_2142_wire(0) /=  '0') else IMC20_1970;
    -- logger for split-operator MUX_2153_inst flow-through 
    process(IMD11_2154) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_2153_inst:flowthrough inputs: " & " BITSEL_u8_u1_2150_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_2150_wire) & " IMC23_1994 = "& Convert_SLV_To_Hex_String(IMC23_1994) & " IMC22_1986 = "& Convert_SLV_To_Hex_String(IMC22_1986) & " outputs:" & " IMD11_2154= "  & Convert_SLV_To_Hex_String(IMD11_2154));
      --
    end process; 
    -- flow-through select operator MUX_2153_inst
    IMD11_2154 <= IMC23_1994 when (BITSEL_u8_u1_2150_wire(0) /=  '0') else IMC22_1986;
    -- logger for split-operator MUX_2161_inst flow-through 
    process(IMD12_2162) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_2161_inst:flowthrough inputs: " & " BITSEL_u8_u1_2158_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_2158_wire) & " IMC25_2010 = "& Convert_SLV_To_Hex_String(IMC25_2010) & " IMC24_2002 = "& Convert_SLV_To_Hex_String(IMC24_2002) & " outputs:" & " IMD12_2162= "  & Convert_SLV_To_Hex_String(IMD12_2162));
      --
    end process; 
    -- flow-through select operator MUX_2161_inst
    IMD12_2162 <= IMC25_2010 when (BITSEL_u8_u1_2158_wire(0) /=  '0') else IMC24_2002;
    -- logger for split-operator MUX_2169_inst flow-through 
    process(IMD13_2170) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_2169_inst:flowthrough inputs: " & " BITSEL_u8_u1_2166_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_2166_wire) & " IMC27_2026 = "& Convert_SLV_To_Hex_String(IMC27_2026) & " IMC26_2018 = "& Convert_SLV_To_Hex_String(IMC26_2018) & " outputs:" & " IMD13_2170= "  & Convert_SLV_To_Hex_String(IMD13_2170));
      --
    end process; 
    -- flow-through select operator MUX_2169_inst
    IMD13_2170 <= IMC27_2026 when (BITSEL_u8_u1_2166_wire(0) /=  '0') else IMC26_2018;
    -- logger for split-operator MUX_2177_inst flow-through 
    process(IMD14_2178) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_2177_inst:flowthrough inputs: " & " BITSEL_u8_u1_2174_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_2174_wire) & " IMC29_2042 = "& Convert_SLV_To_Hex_String(IMC29_2042) & " IMC28_2034 = "& Convert_SLV_To_Hex_String(IMC28_2034) & " outputs:" & " IMD14_2178= "  & Convert_SLV_To_Hex_String(IMD14_2178));
      --
    end process; 
    -- flow-through select operator MUX_2177_inst
    IMD14_2178 <= IMC29_2042 when (BITSEL_u8_u1_2174_wire(0) /=  '0') else IMC28_2034;
    -- logger for split-operator MUX_2185_inst flow-through 
    process(IMD15_2186) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_2185_inst:flowthrough inputs: " & " BITSEL_u8_u1_2182_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_2182_wire) & " IMC31_2058 = "& Convert_SLV_To_Hex_String(IMC31_2058) & " IMC30_2050 = "& Convert_SLV_To_Hex_String(IMC30_2050) & " outputs:" & " IMD15_2186= "  & Convert_SLV_To_Hex_String(IMD15_2186));
      --
    end process; 
    -- flow-through select operator MUX_2185_inst
    IMD15_2186 <= IMC31_2058 when (BITSEL_u8_u1_2182_wire(0) /=  '0') else IMC30_2050;
    -- logger for split-operator MUX_2193_inst flow-through 
    process(IME0_2194) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_2193_inst:flowthrough inputs: " & " BITSEL_u8_u1_2190_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_2190_wire) & " IMD1_2074 = "& Convert_SLV_To_Hex_String(IMD1_2074) & " IMD0_2066 = "& Convert_SLV_To_Hex_String(IMD0_2066) & " outputs:" & " IME0_2194= "  & Convert_SLV_To_Hex_String(IME0_2194));
      --
    end process; 
    -- flow-through select operator MUX_2193_inst
    IME0_2194 <= IMD1_2074 when (BITSEL_u8_u1_2190_wire(0) /=  '0') else IMD0_2066;
    -- logger for split-operator MUX_219_inst flow-through 
    process(IMA20_220) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_219_inst:flowthrough inputs: " & " BITSEL_u8_u1_214_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_214_wire) & " type_cast_216_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_216_wire_constant) & " type_cast_218_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_218_wire_constant) & " outputs:" & " IMA20_220= "  & Convert_SLV_To_Hex_String(IMA20_220));
      --
    end process; 
    -- flow-through select operator MUX_219_inst
    IMA20_220 <= type_cast_216_wire_constant when (BITSEL_u8_u1_214_wire(0) /=  '0') else type_cast_218_wire_constant;
    -- logger for split-operator MUX_2201_inst flow-through 
    process(IME1_2202) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_2201_inst:flowthrough inputs: " & " BITSEL_u8_u1_2198_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_2198_wire) & " IMD3_2090 = "& Convert_SLV_To_Hex_String(IMD3_2090) & " IMD2_2082 = "& Convert_SLV_To_Hex_String(IMD2_2082) & " outputs:" & " IME1_2202= "  & Convert_SLV_To_Hex_String(IME1_2202));
      --
    end process; 
    -- flow-through select operator MUX_2201_inst
    IME1_2202 <= IMD3_2090 when (BITSEL_u8_u1_2198_wire(0) /=  '0') else IMD2_2082;
    -- logger for split-operator MUX_2209_inst flow-through 
    process(IME2_2210) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_2209_inst:flowthrough inputs: " & " BITSEL_u8_u1_2206_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_2206_wire) & " IMD5_2106 = "& Convert_SLV_To_Hex_String(IMD5_2106) & " IMD4_2098 = "& Convert_SLV_To_Hex_String(IMD4_2098) & " outputs:" & " IME2_2210= "  & Convert_SLV_To_Hex_String(IME2_2210));
      --
    end process; 
    -- flow-through select operator MUX_2209_inst
    IME2_2210 <= IMD5_2106 when (BITSEL_u8_u1_2206_wire(0) /=  '0') else IMD4_2098;
    -- logger for split-operator MUX_2217_inst flow-through 
    process(IME3_2218) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_2217_inst:flowthrough inputs: " & " BITSEL_u8_u1_2214_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_2214_wire) & " IMD7_2122 = "& Convert_SLV_To_Hex_String(IMD7_2122) & " IMD6_2114 = "& Convert_SLV_To_Hex_String(IMD6_2114) & " outputs:" & " IME3_2218= "  & Convert_SLV_To_Hex_String(IME3_2218));
      --
    end process; 
    -- flow-through select operator MUX_2217_inst
    IME3_2218 <= IMD7_2122 when (BITSEL_u8_u1_2214_wire(0) /=  '0') else IMD6_2114;
    -- logger for split-operator MUX_2225_inst flow-through 
    process(IME4_2226) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_2225_inst:flowthrough inputs: " & " BITSEL_u8_u1_2222_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_2222_wire) & " IMD9_2138 = "& Convert_SLV_To_Hex_String(IMD9_2138) & " IMD8_2130 = "& Convert_SLV_To_Hex_String(IMD8_2130) & " outputs:" & " IME4_2226= "  & Convert_SLV_To_Hex_String(IME4_2226));
      --
    end process; 
    -- flow-through select operator MUX_2225_inst
    IME4_2226 <= IMD9_2138 when (BITSEL_u8_u1_2222_wire(0) /=  '0') else IMD8_2130;
    -- logger for split-operator MUX_2233_inst flow-through 
    process(IME5_2234) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_2233_inst:flowthrough inputs: " & " BITSEL_u8_u1_2230_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_2230_wire) & " IMD11_2154 = "& Convert_SLV_To_Hex_String(IMD11_2154) & " IMD10_2146 = "& Convert_SLV_To_Hex_String(IMD10_2146) & " outputs:" & " IME5_2234= "  & Convert_SLV_To_Hex_String(IME5_2234));
      --
    end process; 
    -- flow-through select operator MUX_2233_inst
    IME5_2234 <= IMD11_2154 when (BITSEL_u8_u1_2230_wire(0) /=  '0') else IMD10_2146;
    -- logger for split-operator MUX_2241_inst flow-through 
    process(IME6_2242) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_2241_inst:flowthrough inputs: " & " BITSEL_u8_u1_2238_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_2238_wire) & " IMD13_2170 = "& Convert_SLV_To_Hex_String(IMD13_2170) & " IMD12_2162 = "& Convert_SLV_To_Hex_String(IMD12_2162) & " outputs:" & " IME6_2242= "  & Convert_SLV_To_Hex_String(IME6_2242));
      --
    end process; 
    -- flow-through select operator MUX_2241_inst
    IME6_2242 <= IMD13_2170 when (BITSEL_u8_u1_2238_wire(0) /=  '0') else IMD12_2162;
    -- logger for split-operator MUX_2249_inst flow-through 
    process(IME7_2250) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_2249_inst:flowthrough inputs: " & " BITSEL_u8_u1_2246_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_2246_wire) & " IMD15_2186 = "& Convert_SLV_To_Hex_String(IMD15_2186) & " IMD14_2178 = "& Convert_SLV_To_Hex_String(IMD14_2178) & " outputs:" & " IME7_2250= "  & Convert_SLV_To_Hex_String(IME7_2250));
      --
    end process; 
    -- flow-through select operator MUX_2249_inst
    IME7_2250 <= IMD15_2186 when (BITSEL_u8_u1_2246_wire(0) /=  '0') else IMD14_2178;
    -- logger for split-operator MUX_2257_inst flow-through 
    process(IMF0_2258) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_2257_inst:flowthrough inputs: " & " BITSEL_u8_u1_2254_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_2254_wire) & " IME1_2202 = "& Convert_SLV_To_Hex_String(IME1_2202) & " IME0_2194 = "& Convert_SLV_To_Hex_String(IME0_2194) & " outputs:" & " IMF0_2258= "  & Convert_SLV_To_Hex_String(IMF0_2258));
      --
    end process; 
    -- flow-through select operator MUX_2257_inst
    IMF0_2258 <= IME1_2202 when (BITSEL_u8_u1_2254_wire(0) /=  '0') else IME0_2194;
    -- logger for split-operator MUX_2265_inst flow-through 
    process(IMF1_2266) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_2265_inst:flowthrough inputs: " & " BITSEL_u8_u1_2262_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_2262_wire) & " IME3_2218 = "& Convert_SLV_To_Hex_String(IME3_2218) & " IME2_2210 = "& Convert_SLV_To_Hex_String(IME2_2210) & " outputs:" & " IMF1_2266= "  & Convert_SLV_To_Hex_String(IMF1_2266));
      --
    end process; 
    -- flow-through select operator MUX_2265_inst
    IMF1_2266 <= IME3_2218 when (BITSEL_u8_u1_2262_wire(0) /=  '0') else IME2_2210;
    -- logger for split-operator MUX_2273_inst flow-through 
    process(IMF2_2274) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_2273_inst:flowthrough inputs: " & " BITSEL_u8_u1_2270_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_2270_wire) & " IME5_2234 = "& Convert_SLV_To_Hex_String(IME5_2234) & " IME4_2226 = "& Convert_SLV_To_Hex_String(IME4_2226) & " outputs:" & " IMF2_2274= "  & Convert_SLV_To_Hex_String(IMF2_2274));
      --
    end process; 
    -- flow-through select operator MUX_2273_inst
    IMF2_2274 <= IME5_2234 when (BITSEL_u8_u1_2270_wire(0) /=  '0') else IME4_2226;
    -- logger for split-operator MUX_2281_inst flow-through 
    process(IMF3_2282) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_2281_inst:flowthrough inputs: " & " BITSEL_u8_u1_2278_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_2278_wire) & " IME7_2250 = "& Convert_SLV_To_Hex_String(IME7_2250) & " IME6_2242 = "& Convert_SLV_To_Hex_String(IME6_2242) & " outputs:" & " IMF3_2282= "  & Convert_SLV_To_Hex_String(IMF3_2282));
      --
    end process; 
    -- flow-through select operator MUX_2281_inst
    IMF3_2282 <= IME7_2250 when (BITSEL_u8_u1_2278_wire(0) /=  '0') else IME6_2242;
    -- logger for split-operator MUX_2289_inst flow-through 
    process(IMG0_2290) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_2289_inst:flowthrough inputs: " & " BITSEL_u8_u1_2286_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_2286_wire) & " IMF1_2266 = "& Convert_SLV_To_Hex_String(IMF1_2266) & " IMF0_2258 = "& Convert_SLV_To_Hex_String(IMF0_2258) & " outputs:" & " IMG0_2290= "  & Convert_SLV_To_Hex_String(IMG0_2290));
      --
    end process; 
    -- flow-through select operator MUX_2289_inst
    IMG0_2290 <= IMF1_2266 when (BITSEL_u8_u1_2286_wire(0) /=  '0') else IMF0_2258;
    -- logger for split-operator MUX_2297_inst flow-through 
    process(IMG1_2298) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_2297_inst:flowthrough inputs: " & " BITSEL_u8_u1_2294_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_2294_wire) & " IMF3_2282 = "& Convert_SLV_To_Hex_String(IMF3_2282) & " IMF2_2274 = "& Convert_SLV_To_Hex_String(IMF2_2274) & " outputs:" & " IMG1_2298= "  & Convert_SLV_To_Hex_String(IMG1_2298));
      --
    end process; 
    -- flow-through select operator MUX_2297_inst
    IMG1_2298 <= IMF3_2282 when (BITSEL_u8_u1_2294_wire(0) /=  '0') else IMF2_2274;
    -- logger for split-operator MUX_229_inst flow-through 
    process(IMA21_230) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_229_inst:flowthrough inputs: " & " BITSEL_u8_u1_224_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_224_wire) & " type_cast_226_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_226_wire_constant) & " type_cast_228_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_228_wire_constant) & " outputs:" & " IMA21_230= "  & Convert_SLV_To_Hex_String(IMA21_230));
      --
    end process; 
    -- flow-through select operator MUX_229_inst
    IMA21_230 <= type_cast_226_wire_constant when (BITSEL_u8_u1_224_wire(0) /=  '0') else type_cast_228_wire_constant;
    -- logger for split-operator MUX_2305_inst flow-through 
    process(s_out_buffer) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_2305_inst:flowthrough inputs: " & " BITSEL_u8_u1_2302_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_2302_wire) & " IMG1_2298 = "& Convert_SLV_To_Hex_String(IMG1_2298) & " IMG0_2290 = "& Convert_SLV_To_Hex_String(IMG0_2290) & " outputs:" & " s_out_buffer= "  & Convert_SLV_To_Hex_String(s_out_buffer));
      --
    end process; 
    -- flow-through select operator MUX_2305_inst
    s_out_buffer <= IMG1_2298 when (BITSEL_u8_u1_2302_wire(0) /=  '0') else IMG0_2290;
    -- logger for split-operator MUX_239_inst flow-through 
    process(IMA22_240) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_239_inst:flowthrough inputs: " & " BITSEL_u8_u1_234_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_234_wire) & " type_cast_236_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_236_wire_constant) & " type_cast_238_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_238_wire_constant) & " outputs:" & " IMA22_240= "  & Convert_SLV_To_Hex_String(IMA22_240));
      --
    end process; 
    -- flow-through select operator MUX_239_inst
    IMA22_240 <= type_cast_236_wire_constant when (BITSEL_u8_u1_234_wire(0) /=  '0') else type_cast_238_wire_constant;
    -- logger for split-operator MUX_249_inst flow-through 
    process(IMA23_250) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_249_inst:flowthrough inputs: " & " BITSEL_u8_u1_244_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_244_wire) & " type_cast_246_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_246_wire_constant) & " type_cast_248_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_248_wire_constant) & " outputs:" & " IMA23_250= "  & Convert_SLV_To_Hex_String(IMA23_250));
      --
    end process; 
    -- flow-through select operator MUX_249_inst
    IMA23_250 <= type_cast_246_wire_constant when (BITSEL_u8_u1_244_wire(0) /=  '0') else type_cast_248_wire_constant;
    -- logger for split-operator MUX_259_inst flow-through 
    process(IMA24_260) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_259_inst:flowthrough inputs: " & " BITSEL_u8_u1_254_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_254_wire) & " type_cast_256_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_256_wire_constant) & " type_cast_258_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_258_wire_constant) & " outputs:" & " IMA24_260= "  & Convert_SLV_To_Hex_String(IMA24_260));
      --
    end process; 
    -- flow-through select operator MUX_259_inst
    IMA24_260 <= type_cast_256_wire_constant when (BITSEL_u8_u1_254_wire(0) /=  '0') else type_cast_258_wire_constant;
    -- logger for split-operator MUX_269_inst flow-through 
    process(IMA25_270) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_269_inst:flowthrough inputs: " & " BITSEL_u8_u1_264_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_264_wire) & " type_cast_266_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_266_wire_constant) & " type_cast_268_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_268_wire_constant) & " outputs:" & " IMA25_270= "  & Convert_SLV_To_Hex_String(IMA25_270));
      --
    end process; 
    -- flow-through select operator MUX_269_inst
    IMA25_270 <= type_cast_266_wire_constant when (BITSEL_u8_u1_264_wire(0) /=  '0') else type_cast_268_wire_constant;
    -- logger for split-operator MUX_279_inst flow-through 
    process(IMA26_280) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_279_inst:flowthrough inputs: " & " BITSEL_u8_u1_274_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_274_wire) & " type_cast_276_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_276_wire_constant) & " type_cast_278_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_278_wire_constant) & " outputs:" & " IMA26_280= "  & Convert_SLV_To_Hex_String(IMA26_280));
      --
    end process; 
    -- flow-through select operator MUX_279_inst
    IMA26_280 <= type_cast_276_wire_constant when (BITSEL_u8_u1_274_wire(0) /=  '0') else type_cast_278_wire_constant;
    -- logger for split-operator MUX_289_inst flow-through 
    process(IMA27_290) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_289_inst:flowthrough inputs: " & " BITSEL_u8_u1_284_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_284_wire) & " type_cast_286_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_286_wire_constant) & " type_cast_288_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_288_wire_constant) & " outputs:" & " IMA27_290= "  & Convert_SLV_To_Hex_String(IMA27_290));
      --
    end process; 
    -- flow-through select operator MUX_289_inst
    IMA27_290 <= type_cast_286_wire_constant when (BITSEL_u8_u1_284_wire(0) /=  '0') else type_cast_288_wire_constant;
    -- logger for split-operator MUX_299_inst flow-through 
    process(IMA28_300) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_299_inst:flowthrough inputs: " & " BITSEL_u8_u1_294_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_294_wire) & " type_cast_296_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_296_wire_constant) & " type_cast_298_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_298_wire_constant) & " outputs:" & " IMA28_300= "  & Convert_SLV_To_Hex_String(IMA28_300));
      --
    end process; 
    -- flow-through select operator MUX_299_inst
    IMA28_300 <= type_cast_296_wire_constant when (BITSEL_u8_u1_294_wire(0) /=  '0') else type_cast_298_wire_constant;
    -- logger for split-operator MUX_29_inst flow-through 
    process(IMA1_30) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_29_inst:flowthrough inputs: " & " BITSEL_u8_u1_24_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_24_wire) & " type_cast_26_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_26_wire_constant) & " type_cast_28_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_28_wire_constant) & " outputs:" & " IMA1_30= "  & Convert_SLV_To_Hex_String(IMA1_30));
      --
    end process; 
    -- flow-through select operator MUX_29_inst
    IMA1_30 <= type_cast_26_wire_constant when (BITSEL_u8_u1_24_wire(0) /=  '0') else type_cast_28_wire_constant;
    -- logger for split-operator MUX_309_inst flow-through 
    process(IMA29_310) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_309_inst:flowthrough inputs: " & " BITSEL_u8_u1_304_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_304_wire) & " type_cast_306_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_306_wire_constant) & " type_cast_308_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_308_wire_constant) & " outputs:" & " IMA29_310= "  & Convert_SLV_To_Hex_String(IMA29_310));
      --
    end process; 
    -- flow-through select operator MUX_309_inst
    IMA29_310 <= type_cast_306_wire_constant when (BITSEL_u8_u1_304_wire(0) /=  '0') else type_cast_308_wire_constant;
    -- logger for split-operator MUX_319_inst flow-through 
    process(IMA30_320) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_319_inst:flowthrough inputs: " & " BITSEL_u8_u1_314_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_314_wire) & " type_cast_316_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_316_wire_constant) & " type_cast_318_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_318_wire_constant) & " outputs:" & " IMA30_320= "  & Convert_SLV_To_Hex_String(IMA30_320));
      --
    end process; 
    -- flow-through select operator MUX_319_inst
    IMA30_320 <= type_cast_316_wire_constant when (BITSEL_u8_u1_314_wire(0) /=  '0') else type_cast_318_wire_constant;
    -- logger for split-operator MUX_329_inst flow-through 
    process(IMA31_330) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_329_inst:flowthrough inputs: " & " BITSEL_u8_u1_324_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_324_wire) & " type_cast_326_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_326_wire_constant) & " type_cast_328_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_328_wire_constant) & " outputs:" & " IMA31_330= "  & Convert_SLV_To_Hex_String(IMA31_330));
      --
    end process; 
    -- flow-through select operator MUX_329_inst
    IMA31_330 <= type_cast_326_wire_constant when (BITSEL_u8_u1_324_wire(0) /=  '0') else type_cast_328_wire_constant;
    -- logger for split-operator MUX_339_inst flow-through 
    process(IMA32_340) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_339_inst:flowthrough inputs: " & " BITSEL_u8_u1_334_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_334_wire) & " type_cast_336_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_336_wire_constant) & " type_cast_338_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_338_wire_constant) & " outputs:" & " IMA32_340= "  & Convert_SLV_To_Hex_String(IMA32_340));
      --
    end process; 
    -- flow-through select operator MUX_339_inst
    IMA32_340 <= type_cast_336_wire_constant when (BITSEL_u8_u1_334_wire(0) /=  '0') else type_cast_338_wire_constant;
    -- logger for split-operator MUX_349_inst flow-through 
    process(IMA33_350) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_349_inst:flowthrough inputs: " & " BITSEL_u8_u1_344_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_344_wire) & " type_cast_346_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_346_wire_constant) & " type_cast_348_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_348_wire_constant) & " outputs:" & " IMA33_350= "  & Convert_SLV_To_Hex_String(IMA33_350));
      --
    end process; 
    -- flow-through select operator MUX_349_inst
    IMA33_350 <= type_cast_346_wire_constant when (BITSEL_u8_u1_344_wire(0) /=  '0') else type_cast_348_wire_constant;
    -- logger for split-operator MUX_359_inst flow-through 
    process(IMA34_360) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_359_inst:flowthrough inputs: " & " BITSEL_u8_u1_354_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_354_wire) & " type_cast_356_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_356_wire_constant) & " type_cast_358_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_358_wire_constant) & " outputs:" & " IMA34_360= "  & Convert_SLV_To_Hex_String(IMA34_360));
      --
    end process; 
    -- flow-through select operator MUX_359_inst
    IMA34_360 <= type_cast_356_wire_constant when (BITSEL_u8_u1_354_wire(0) /=  '0') else type_cast_358_wire_constant;
    -- logger for split-operator MUX_369_inst flow-through 
    process(IMA35_370) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_369_inst:flowthrough inputs: " & " BITSEL_u8_u1_364_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_364_wire) & " type_cast_366_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_366_wire_constant) & " type_cast_368_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_368_wire_constant) & " outputs:" & " IMA35_370= "  & Convert_SLV_To_Hex_String(IMA35_370));
      --
    end process; 
    -- flow-through select operator MUX_369_inst
    IMA35_370 <= type_cast_366_wire_constant when (BITSEL_u8_u1_364_wire(0) /=  '0') else type_cast_368_wire_constant;
    -- logger for split-operator MUX_379_inst flow-through 
    process(IMA36_380) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_379_inst:flowthrough inputs: " & " BITSEL_u8_u1_374_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_374_wire) & " type_cast_376_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_376_wire_constant) & " type_cast_378_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_378_wire_constant) & " outputs:" & " IMA36_380= "  & Convert_SLV_To_Hex_String(IMA36_380));
      --
    end process; 
    -- flow-through select operator MUX_379_inst
    IMA36_380 <= type_cast_376_wire_constant when (BITSEL_u8_u1_374_wire(0) /=  '0') else type_cast_378_wire_constant;
    -- logger for split-operator MUX_389_inst flow-through 
    process(IMA37_390) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_389_inst:flowthrough inputs: " & " BITSEL_u8_u1_384_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_384_wire) & " type_cast_386_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_386_wire_constant) & " type_cast_388_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_388_wire_constant) & " outputs:" & " IMA37_390= "  & Convert_SLV_To_Hex_String(IMA37_390));
      --
    end process; 
    -- flow-through select operator MUX_389_inst
    IMA37_390 <= type_cast_386_wire_constant when (BITSEL_u8_u1_384_wire(0) /=  '0') else type_cast_388_wire_constant;
    -- logger for split-operator MUX_399_inst flow-through 
    process(IMA38_400) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_399_inst:flowthrough inputs: " & " BITSEL_u8_u1_394_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_394_wire) & " type_cast_396_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_396_wire_constant) & " type_cast_398_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_398_wire_constant) & " outputs:" & " IMA38_400= "  & Convert_SLV_To_Hex_String(IMA38_400));
      --
    end process; 
    -- flow-through select operator MUX_399_inst
    IMA38_400 <= type_cast_396_wire_constant when (BITSEL_u8_u1_394_wire(0) /=  '0') else type_cast_398_wire_constant;
    -- logger for split-operator MUX_39_inst flow-through 
    process(IMA2_40) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_39_inst:flowthrough inputs: " & " BITSEL_u8_u1_34_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_34_wire) & " type_cast_36_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_36_wire_constant) & " type_cast_38_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_38_wire_constant) & " outputs:" & " IMA2_40= "  & Convert_SLV_To_Hex_String(IMA2_40));
      --
    end process; 
    -- flow-through select operator MUX_39_inst
    IMA2_40 <= type_cast_36_wire_constant when (BITSEL_u8_u1_34_wire(0) /=  '0') else type_cast_38_wire_constant;
    -- logger for split-operator MUX_409_inst flow-through 
    process(IMA39_410) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_409_inst:flowthrough inputs: " & " BITSEL_u8_u1_404_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_404_wire) & " type_cast_406_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_406_wire_constant) & " type_cast_408_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_408_wire_constant) & " outputs:" & " IMA39_410= "  & Convert_SLV_To_Hex_String(IMA39_410));
      --
    end process; 
    -- flow-through select operator MUX_409_inst
    IMA39_410 <= type_cast_406_wire_constant when (BITSEL_u8_u1_404_wire(0) /=  '0') else type_cast_408_wire_constant;
    -- logger for split-operator MUX_419_inst flow-through 
    process(IMA40_420) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_419_inst:flowthrough inputs: " & " BITSEL_u8_u1_414_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_414_wire) & " type_cast_416_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_416_wire_constant) & " type_cast_418_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_418_wire_constant) & " outputs:" & " IMA40_420= "  & Convert_SLV_To_Hex_String(IMA40_420));
      --
    end process; 
    -- flow-through select operator MUX_419_inst
    IMA40_420 <= type_cast_416_wire_constant when (BITSEL_u8_u1_414_wire(0) /=  '0') else type_cast_418_wire_constant;
    -- logger for split-operator MUX_429_inst flow-through 
    process(IMA41_430) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_429_inst:flowthrough inputs: " & " BITSEL_u8_u1_424_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_424_wire) & " type_cast_426_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_426_wire_constant) & " type_cast_428_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_428_wire_constant) & " outputs:" & " IMA41_430= "  & Convert_SLV_To_Hex_String(IMA41_430));
      --
    end process; 
    -- flow-through select operator MUX_429_inst
    IMA41_430 <= type_cast_426_wire_constant when (BITSEL_u8_u1_424_wire(0) /=  '0') else type_cast_428_wire_constant;
    -- logger for split-operator MUX_439_inst flow-through 
    process(IMA42_440) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_439_inst:flowthrough inputs: " & " BITSEL_u8_u1_434_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_434_wire) & " type_cast_436_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_436_wire_constant) & " type_cast_438_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_438_wire_constant) & " outputs:" & " IMA42_440= "  & Convert_SLV_To_Hex_String(IMA42_440));
      --
    end process; 
    -- flow-through select operator MUX_439_inst
    IMA42_440 <= type_cast_436_wire_constant when (BITSEL_u8_u1_434_wire(0) /=  '0') else type_cast_438_wire_constant;
    -- logger for split-operator MUX_449_inst flow-through 
    process(IMA43_450) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_449_inst:flowthrough inputs: " & " BITSEL_u8_u1_444_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_444_wire) & " type_cast_446_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_446_wire_constant) & " type_cast_448_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_448_wire_constant) & " outputs:" & " IMA43_450= "  & Convert_SLV_To_Hex_String(IMA43_450));
      --
    end process; 
    -- flow-through select operator MUX_449_inst
    IMA43_450 <= type_cast_446_wire_constant when (BITSEL_u8_u1_444_wire(0) /=  '0') else type_cast_448_wire_constant;
    -- logger for split-operator MUX_459_inst flow-through 
    process(IMA44_460) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_459_inst:flowthrough inputs: " & " BITSEL_u8_u1_454_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_454_wire) & " type_cast_456_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_456_wire_constant) & " type_cast_458_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_458_wire_constant) & " outputs:" & " IMA44_460= "  & Convert_SLV_To_Hex_String(IMA44_460));
      --
    end process; 
    -- flow-through select operator MUX_459_inst
    IMA44_460 <= type_cast_456_wire_constant when (BITSEL_u8_u1_454_wire(0) /=  '0') else type_cast_458_wire_constant;
    -- logger for split-operator MUX_469_inst flow-through 
    process(IMA45_470) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_469_inst:flowthrough inputs: " & " BITSEL_u8_u1_464_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_464_wire) & " type_cast_466_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_466_wire_constant) & " type_cast_468_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_468_wire_constant) & " outputs:" & " IMA45_470= "  & Convert_SLV_To_Hex_String(IMA45_470));
      --
    end process; 
    -- flow-through select operator MUX_469_inst
    IMA45_470 <= type_cast_466_wire_constant when (BITSEL_u8_u1_464_wire(0) /=  '0') else type_cast_468_wire_constant;
    -- logger for split-operator MUX_479_inst flow-through 
    process(IMA46_480) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_479_inst:flowthrough inputs: " & " BITSEL_u8_u1_474_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_474_wire) & " type_cast_476_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_476_wire_constant) & " type_cast_478_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_478_wire_constant) & " outputs:" & " IMA46_480= "  & Convert_SLV_To_Hex_String(IMA46_480));
      --
    end process; 
    -- flow-through select operator MUX_479_inst
    IMA46_480 <= type_cast_476_wire_constant when (BITSEL_u8_u1_474_wire(0) /=  '0') else type_cast_478_wire_constant;
    -- logger for split-operator MUX_489_inst flow-through 
    process(IMA47_490) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_489_inst:flowthrough inputs: " & " BITSEL_u8_u1_484_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_484_wire) & " type_cast_486_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_486_wire_constant) & " type_cast_488_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_488_wire_constant) & " outputs:" & " IMA47_490= "  & Convert_SLV_To_Hex_String(IMA47_490));
      --
    end process; 
    -- flow-through select operator MUX_489_inst
    IMA47_490 <= type_cast_486_wire_constant when (BITSEL_u8_u1_484_wire(0) /=  '0') else type_cast_488_wire_constant;
    -- logger for split-operator MUX_499_inst flow-through 
    process(IMA48_500) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_499_inst:flowthrough inputs: " & " BITSEL_u8_u1_494_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_494_wire) & " type_cast_496_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_496_wire_constant) & " type_cast_498_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_498_wire_constant) & " outputs:" & " IMA48_500= "  & Convert_SLV_To_Hex_String(IMA48_500));
      --
    end process; 
    -- flow-through select operator MUX_499_inst
    IMA48_500 <= type_cast_496_wire_constant when (BITSEL_u8_u1_494_wire(0) /=  '0') else type_cast_498_wire_constant;
    -- logger for split-operator MUX_49_inst flow-through 
    process(IMA3_50) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_49_inst:flowthrough inputs: " & " BITSEL_u8_u1_44_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_44_wire) & " type_cast_46_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_46_wire_constant) & " type_cast_48_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_48_wire_constant) & " outputs:" & " IMA3_50= "  & Convert_SLV_To_Hex_String(IMA3_50));
      --
    end process; 
    -- flow-through select operator MUX_49_inst
    IMA3_50 <= type_cast_46_wire_constant when (BITSEL_u8_u1_44_wire(0) /=  '0') else type_cast_48_wire_constant;
    -- logger for split-operator MUX_509_inst flow-through 
    process(IMA49_510) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_509_inst:flowthrough inputs: " & " BITSEL_u8_u1_504_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_504_wire) & " type_cast_506_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_506_wire_constant) & " type_cast_508_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_508_wire_constant) & " outputs:" & " IMA49_510= "  & Convert_SLV_To_Hex_String(IMA49_510));
      --
    end process; 
    -- flow-through select operator MUX_509_inst
    IMA49_510 <= type_cast_506_wire_constant when (BITSEL_u8_u1_504_wire(0) /=  '0') else type_cast_508_wire_constant;
    -- logger for split-operator MUX_519_inst flow-through 
    process(IMA50_520) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_519_inst:flowthrough inputs: " & " BITSEL_u8_u1_514_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_514_wire) & " type_cast_516_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_516_wire_constant) & " type_cast_518_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_518_wire_constant) & " outputs:" & " IMA50_520= "  & Convert_SLV_To_Hex_String(IMA50_520));
      --
    end process; 
    -- flow-through select operator MUX_519_inst
    IMA50_520 <= type_cast_516_wire_constant when (BITSEL_u8_u1_514_wire(0) /=  '0') else type_cast_518_wire_constant;
    -- logger for split-operator MUX_529_inst flow-through 
    process(IMA51_530) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_529_inst:flowthrough inputs: " & " BITSEL_u8_u1_524_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_524_wire) & " type_cast_526_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_526_wire_constant) & " type_cast_528_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_528_wire_constant) & " outputs:" & " IMA51_530= "  & Convert_SLV_To_Hex_String(IMA51_530));
      --
    end process; 
    -- flow-through select operator MUX_529_inst
    IMA51_530 <= type_cast_526_wire_constant when (BITSEL_u8_u1_524_wire(0) /=  '0') else type_cast_528_wire_constant;
    -- logger for split-operator MUX_539_inst flow-through 
    process(IMA52_540) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_539_inst:flowthrough inputs: " & " BITSEL_u8_u1_534_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_534_wire) & " type_cast_536_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_536_wire_constant) & " type_cast_538_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_538_wire_constant) & " outputs:" & " IMA52_540= "  & Convert_SLV_To_Hex_String(IMA52_540));
      --
    end process; 
    -- flow-through select operator MUX_539_inst
    IMA52_540 <= type_cast_536_wire_constant when (BITSEL_u8_u1_534_wire(0) /=  '0') else type_cast_538_wire_constant;
    -- logger for split-operator MUX_549_inst flow-through 
    process(IMA53_550) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_549_inst:flowthrough inputs: " & " BITSEL_u8_u1_544_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_544_wire) & " type_cast_546_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_546_wire_constant) & " type_cast_548_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_548_wire_constant) & " outputs:" & " IMA53_550= "  & Convert_SLV_To_Hex_String(IMA53_550));
      --
    end process; 
    -- flow-through select operator MUX_549_inst
    IMA53_550 <= type_cast_546_wire_constant when (BITSEL_u8_u1_544_wire(0) /=  '0') else type_cast_548_wire_constant;
    -- logger for split-operator MUX_559_inst flow-through 
    process(IMA54_560) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_559_inst:flowthrough inputs: " & " BITSEL_u8_u1_554_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_554_wire) & " type_cast_556_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_556_wire_constant) & " type_cast_558_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_558_wire_constant) & " outputs:" & " IMA54_560= "  & Convert_SLV_To_Hex_String(IMA54_560));
      --
    end process; 
    -- flow-through select operator MUX_559_inst
    IMA54_560 <= type_cast_556_wire_constant when (BITSEL_u8_u1_554_wire(0) /=  '0') else type_cast_558_wire_constant;
    -- logger for split-operator MUX_569_inst flow-through 
    process(IMA55_570) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_569_inst:flowthrough inputs: " & " BITSEL_u8_u1_564_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_564_wire) & " type_cast_566_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_566_wire_constant) & " type_cast_568_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_568_wire_constant) & " outputs:" & " IMA55_570= "  & Convert_SLV_To_Hex_String(IMA55_570));
      --
    end process; 
    -- flow-through select operator MUX_569_inst
    IMA55_570 <= type_cast_566_wire_constant when (BITSEL_u8_u1_564_wire(0) /=  '0') else type_cast_568_wire_constant;
    -- logger for split-operator MUX_579_inst flow-through 
    process(IMA56_580) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_579_inst:flowthrough inputs: " & " BITSEL_u8_u1_574_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_574_wire) & " type_cast_576_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_576_wire_constant) & " type_cast_578_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_578_wire_constant) & " outputs:" & " IMA56_580= "  & Convert_SLV_To_Hex_String(IMA56_580));
      --
    end process; 
    -- flow-through select operator MUX_579_inst
    IMA56_580 <= type_cast_576_wire_constant when (BITSEL_u8_u1_574_wire(0) /=  '0') else type_cast_578_wire_constant;
    -- logger for split-operator MUX_589_inst flow-through 
    process(IMA57_590) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_589_inst:flowthrough inputs: " & " BITSEL_u8_u1_584_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_584_wire) & " type_cast_586_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_586_wire_constant) & " type_cast_588_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_588_wire_constant) & " outputs:" & " IMA57_590= "  & Convert_SLV_To_Hex_String(IMA57_590));
      --
    end process; 
    -- flow-through select operator MUX_589_inst
    IMA57_590 <= type_cast_586_wire_constant when (BITSEL_u8_u1_584_wire(0) /=  '0') else type_cast_588_wire_constant;
    -- logger for split-operator MUX_599_inst flow-through 
    process(IMA58_600) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_599_inst:flowthrough inputs: " & " BITSEL_u8_u1_594_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_594_wire) & " type_cast_596_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_596_wire_constant) & " type_cast_598_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_598_wire_constant) & " outputs:" & " IMA58_600= "  & Convert_SLV_To_Hex_String(IMA58_600));
      --
    end process; 
    -- flow-through select operator MUX_599_inst
    IMA58_600 <= type_cast_596_wire_constant when (BITSEL_u8_u1_594_wire(0) /=  '0') else type_cast_598_wire_constant;
    -- logger for split-operator MUX_59_inst flow-through 
    process(IMA4_60) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_59_inst:flowthrough inputs: " & " BITSEL_u8_u1_54_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_54_wire) & " type_cast_56_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_56_wire_constant) & " type_cast_58_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_58_wire_constant) & " outputs:" & " IMA4_60= "  & Convert_SLV_To_Hex_String(IMA4_60));
      --
    end process; 
    -- flow-through select operator MUX_59_inst
    IMA4_60 <= type_cast_56_wire_constant when (BITSEL_u8_u1_54_wire(0) /=  '0') else type_cast_58_wire_constant;
    -- logger for split-operator MUX_609_inst flow-through 
    process(IMA59_610) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_609_inst:flowthrough inputs: " & " BITSEL_u8_u1_604_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_604_wire) & " type_cast_606_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_606_wire_constant) & " type_cast_608_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_608_wire_constant) & " outputs:" & " IMA59_610= "  & Convert_SLV_To_Hex_String(IMA59_610));
      --
    end process; 
    -- flow-through select operator MUX_609_inst
    IMA59_610 <= type_cast_606_wire_constant when (BITSEL_u8_u1_604_wire(0) /=  '0') else type_cast_608_wire_constant;
    -- logger for split-operator MUX_619_inst flow-through 
    process(IMA60_620) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_619_inst:flowthrough inputs: " & " BITSEL_u8_u1_614_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_614_wire) & " type_cast_616_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_616_wire_constant) & " type_cast_618_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_618_wire_constant) & " outputs:" & " IMA60_620= "  & Convert_SLV_To_Hex_String(IMA60_620));
      --
    end process; 
    -- flow-through select operator MUX_619_inst
    IMA60_620 <= type_cast_616_wire_constant when (BITSEL_u8_u1_614_wire(0) /=  '0') else type_cast_618_wire_constant;
    -- logger for split-operator MUX_629_inst flow-through 
    process(IMA61_630) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_629_inst:flowthrough inputs: " & " BITSEL_u8_u1_624_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_624_wire) & " type_cast_626_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_626_wire_constant) & " type_cast_628_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_628_wire_constant) & " outputs:" & " IMA61_630= "  & Convert_SLV_To_Hex_String(IMA61_630));
      --
    end process; 
    -- flow-through select operator MUX_629_inst
    IMA61_630 <= type_cast_626_wire_constant when (BITSEL_u8_u1_624_wire(0) /=  '0') else type_cast_628_wire_constant;
    -- logger for split-operator MUX_639_inst flow-through 
    process(IMA62_640) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_639_inst:flowthrough inputs: " & " BITSEL_u8_u1_634_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_634_wire) & " type_cast_636_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_636_wire_constant) & " type_cast_638_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_638_wire_constant) & " outputs:" & " IMA62_640= "  & Convert_SLV_To_Hex_String(IMA62_640));
      --
    end process; 
    -- flow-through select operator MUX_639_inst
    IMA62_640 <= type_cast_636_wire_constant when (BITSEL_u8_u1_634_wire(0) /=  '0') else type_cast_638_wire_constant;
    -- logger for split-operator MUX_649_inst flow-through 
    process(IMA63_650) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_649_inst:flowthrough inputs: " & " BITSEL_u8_u1_644_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_644_wire) & " type_cast_646_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_646_wire_constant) & " type_cast_648_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_648_wire_constant) & " outputs:" & " IMA63_650= "  & Convert_SLV_To_Hex_String(IMA63_650));
      --
    end process; 
    -- flow-through select operator MUX_649_inst
    IMA63_650 <= type_cast_646_wire_constant when (BITSEL_u8_u1_644_wire(0) /=  '0') else type_cast_648_wire_constant;
    -- logger for split-operator MUX_659_inst flow-through 
    process(IMA64_660) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_659_inst:flowthrough inputs: " & " BITSEL_u8_u1_654_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_654_wire) & " type_cast_656_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_656_wire_constant) & " type_cast_658_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_658_wire_constant) & " outputs:" & " IMA64_660= "  & Convert_SLV_To_Hex_String(IMA64_660));
      --
    end process; 
    -- flow-through select operator MUX_659_inst
    IMA64_660 <= type_cast_656_wire_constant when (BITSEL_u8_u1_654_wire(0) /=  '0') else type_cast_658_wire_constant;
    -- logger for split-operator MUX_669_inst flow-through 
    process(IMA65_670) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_669_inst:flowthrough inputs: " & " BITSEL_u8_u1_664_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_664_wire) & " type_cast_666_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_666_wire_constant) & " type_cast_668_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_668_wire_constant) & " outputs:" & " IMA65_670= "  & Convert_SLV_To_Hex_String(IMA65_670));
      --
    end process; 
    -- flow-through select operator MUX_669_inst
    IMA65_670 <= type_cast_666_wire_constant when (BITSEL_u8_u1_664_wire(0) /=  '0') else type_cast_668_wire_constant;
    -- logger for split-operator MUX_679_inst flow-through 
    process(IMA66_680) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_679_inst:flowthrough inputs: " & " BITSEL_u8_u1_674_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_674_wire) & " type_cast_676_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_676_wire_constant) & " type_cast_678_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_678_wire_constant) & " outputs:" & " IMA66_680= "  & Convert_SLV_To_Hex_String(IMA66_680));
      --
    end process; 
    -- flow-through select operator MUX_679_inst
    IMA66_680 <= type_cast_676_wire_constant when (BITSEL_u8_u1_674_wire(0) /=  '0') else type_cast_678_wire_constant;
    -- logger for split-operator MUX_689_inst flow-through 
    process(IMA67_690) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_689_inst:flowthrough inputs: " & " BITSEL_u8_u1_684_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_684_wire) & " type_cast_686_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_686_wire_constant) & " type_cast_688_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_688_wire_constant) & " outputs:" & " IMA67_690= "  & Convert_SLV_To_Hex_String(IMA67_690));
      --
    end process; 
    -- flow-through select operator MUX_689_inst
    IMA67_690 <= type_cast_686_wire_constant when (BITSEL_u8_u1_684_wire(0) /=  '0') else type_cast_688_wire_constant;
    -- logger for split-operator MUX_699_inst flow-through 
    process(IMA68_700) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_699_inst:flowthrough inputs: " & " BITSEL_u8_u1_694_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_694_wire) & " type_cast_696_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_696_wire_constant) & " type_cast_698_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_698_wire_constant) & " outputs:" & " IMA68_700= "  & Convert_SLV_To_Hex_String(IMA68_700));
      --
    end process; 
    -- flow-through select operator MUX_699_inst
    IMA68_700 <= type_cast_696_wire_constant when (BITSEL_u8_u1_694_wire(0) /=  '0') else type_cast_698_wire_constant;
    -- logger for split-operator MUX_69_inst flow-through 
    process(IMA5_70) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_69_inst:flowthrough inputs: " & " BITSEL_u8_u1_64_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_64_wire) & " type_cast_66_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_66_wire_constant) & " type_cast_68_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_68_wire_constant) & " outputs:" & " IMA5_70= "  & Convert_SLV_To_Hex_String(IMA5_70));
      --
    end process; 
    -- flow-through select operator MUX_69_inst
    IMA5_70 <= type_cast_66_wire_constant when (BITSEL_u8_u1_64_wire(0) /=  '0') else type_cast_68_wire_constant;
    -- logger for split-operator MUX_709_inst flow-through 
    process(IMA69_710) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_709_inst:flowthrough inputs: " & " BITSEL_u8_u1_704_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_704_wire) & " type_cast_706_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_706_wire_constant) & " type_cast_708_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_708_wire_constant) & " outputs:" & " IMA69_710= "  & Convert_SLV_To_Hex_String(IMA69_710));
      --
    end process; 
    -- flow-through select operator MUX_709_inst
    IMA69_710 <= type_cast_706_wire_constant when (BITSEL_u8_u1_704_wire(0) /=  '0') else type_cast_708_wire_constant;
    -- logger for split-operator MUX_719_inst flow-through 
    process(IMA70_720) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_719_inst:flowthrough inputs: " & " BITSEL_u8_u1_714_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_714_wire) & " type_cast_716_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_716_wire_constant) & " type_cast_718_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_718_wire_constant) & " outputs:" & " IMA70_720= "  & Convert_SLV_To_Hex_String(IMA70_720));
      --
    end process; 
    -- flow-through select operator MUX_719_inst
    IMA70_720 <= type_cast_716_wire_constant when (BITSEL_u8_u1_714_wire(0) /=  '0') else type_cast_718_wire_constant;
    -- logger for split-operator MUX_729_inst flow-through 
    process(IMA71_730) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_729_inst:flowthrough inputs: " & " BITSEL_u8_u1_724_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_724_wire) & " type_cast_726_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_726_wire_constant) & " type_cast_728_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_728_wire_constant) & " outputs:" & " IMA71_730= "  & Convert_SLV_To_Hex_String(IMA71_730));
      --
    end process; 
    -- flow-through select operator MUX_729_inst
    IMA71_730 <= type_cast_726_wire_constant when (BITSEL_u8_u1_724_wire(0) /=  '0') else type_cast_728_wire_constant;
    -- logger for split-operator MUX_739_inst flow-through 
    process(IMA72_740) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_739_inst:flowthrough inputs: " & " BITSEL_u8_u1_734_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_734_wire) & " type_cast_736_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_736_wire_constant) & " type_cast_738_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_738_wire_constant) & " outputs:" & " IMA72_740= "  & Convert_SLV_To_Hex_String(IMA72_740));
      --
    end process; 
    -- flow-through select operator MUX_739_inst
    IMA72_740 <= type_cast_736_wire_constant when (BITSEL_u8_u1_734_wire(0) /=  '0') else type_cast_738_wire_constant;
    -- logger for split-operator MUX_749_inst flow-through 
    process(IMA73_750) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_749_inst:flowthrough inputs: " & " BITSEL_u8_u1_744_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_744_wire) & " type_cast_746_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_746_wire_constant) & " type_cast_748_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_748_wire_constant) & " outputs:" & " IMA73_750= "  & Convert_SLV_To_Hex_String(IMA73_750));
      --
    end process; 
    -- flow-through select operator MUX_749_inst
    IMA73_750 <= type_cast_746_wire_constant when (BITSEL_u8_u1_744_wire(0) /=  '0') else type_cast_748_wire_constant;
    -- logger for split-operator MUX_759_inst flow-through 
    process(IMA74_760) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_759_inst:flowthrough inputs: " & " BITSEL_u8_u1_754_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_754_wire) & " type_cast_756_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_756_wire_constant) & " type_cast_758_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_758_wire_constant) & " outputs:" & " IMA74_760= "  & Convert_SLV_To_Hex_String(IMA74_760));
      --
    end process; 
    -- flow-through select operator MUX_759_inst
    IMA74_760 <= type_cast_756_wire_constant when (BITSEL_u8_u1_754_wire(0) /=  '0') else type_cast_758_wire_constant;
    -- logger for split-operator MUX_769_inst flow-through 
    process(IMA75_770) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_769_inst:flowthrough inputs: " & " BITSEL_u8_u1_764_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_764_wire) & " type_cast_766_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_766_wire_constant) & " type_cast_768_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_768_wire_constant) & " outputs:" & " IMA75_770= "  & Convert_SLV_To_Hex_String(IMA75_770));
      --
    end process; 
    -- flow-through select operator MUX_769_inst
    IMA75_770 <= type_cast_766_wire_constant when (BITSEL_u8_u1_764_wire(0) /=  '0') else type_cast_768_wire_constant;
    -- logger for split-operator MUX_779_inst flow-through 
    process(IMA76_780) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_779_inst:flowthrough inputs: " & " BITSEL_u8_u1_774_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_774_wire) & " type_cast_776_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_776_wire_constant) & " type_cast_778_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_778_wire_constant) & " outputs:" & " IMA76_780= "  & Convert_SLV_To_Hex_String(IMA76_780));
      --
    end process; 
    -- flow-through select operator MUX_779_inst
    IMA76_780 <= type_cast_776_wire_constant when (BITSEL_u8_u1_774_wire(0) /=  '0') else type_cast_778_wire_constant;
    -- logger for split-operator MUX_789_inst flow-through 
    process(IMA77_790) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_789_inst:flowthrough inputs: " & " BITSEL_u8_u1_784_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_784_wire) & " type_cast_786_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_786_wire_constant) & " type_cast_788_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_788_wire_constant) & " outputs:" & " IMA77_790= "  & Convert_SLV_To_Hex_String(IMA77_790));
      --
    end process; 
    -- flow-through select operator MUX_789_inst
    IMA77_790 <= type_cast_786_wire_constant when (BITSEL_u8_u1_784_wire(0) /=  '0') else type_cast_788_wire_constant;
    -- logger for split-operator MUX_799_inst flow-through 
    process(IMA78_800) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_799_inst:flowthrough inputs: " & " BITSEL_u8_u1_794_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_794_wire) & " type_cast_796_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_796_wire_constant) & " type_cast_798_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_798_wire_constant) & " outputs:" & " IMA78_800= "  & Convert_SLV_To_Hex_String(IMA78_800));
      --
    end process; 
    -- flow-through select operator MUX_799_inst
    IMA78_800 <= type_cast_796_wire_constant when (BITSEL_u8_u1_794_wire(0) /=  '0') else type_cast_798_wire_constant;
    -- logger for split-operator MUX_79_inst flow-through 
    process(IMA6_80) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_79_inst:flowthrough inputs: " & " BITSEL_u8_u1_74_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_74_wire) & " type_cast_76_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_76_wire_constant) & " type_cast_78_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_78_wire_constant) & " outputs:" & " IMA6_80= "  & Convert_SLV_To_Hex_String(IMA6_80));
      --
    end process; 
    -- flow-through select operator MUX_79_inst
    IMA6_80 <= type_cast_76_wire_constant when (BITSEL_u8_u1_74_wire(0) /=  '0') else type_cast_78_wire_constant;
    -- logger for split-operator MUX_809_inst flow-through 
    process(IMA79_810) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_809_inst:flowthrough inputs: " & " BITSEL_u8_u1_804_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_804_wire) & " type_cast_806_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_806_wire_constant) & " type_cast_808_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_808_wire_constant) & " outputs:" & " IMA79_810= "  & Convert_SLV_To_Hex_String(IMA79_810));
      --
    end process; 
    -- flow-through select operator MUX_809_inst
    IMA79_810 <= type_cast_806_wire_constant when (BITSEL_u8_u1_804_wire(0) /=  '0') else type_cast_808_wire_constant;
    -- logger for split-operator MUX_819_inst flow-through 
    process(IMA80_820) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_819_inst:flowthrough inputs: " & " BITSEL_u8_u1_814_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_814_wire) & " type_cast_816_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_816_wire_constant) & " type_cast_818_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_818_wire_constant) & " outputs:" & " IMA80_820= "  & Convert_SLV_To_Hex_String(IMA80_820));
      --
    end process; 
    -- flow-through select operator MUX_819_inst
    IMA80_820 <= type_cast_816_wire_constant when (BITSEL_u8_u1_814_wire(0) /=  '0') else type_cast_818_wire_constant;
    -- logger for split-operator MUX_829_inst flow-through 
    process(IMA81_830) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_829_inst:flowthrough inputs: " & " BITSEL_u8_u1_824_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_824_wire) & " type_cast_826_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_826_wire_constant) & " type_cast_828_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_828_wire_constant) & " outputs:" & " IMA81_830= "  & Convert_SLV_To_Hex_String(IMA81_830));
      --
    end process; 
    -- flow-through select operator MUX_829_inst
    IMA81_830 <= type_cast_826_wire_constant when (BITSEL_u8_u1_824_wire(0) /=  '0') else type_cast_828_wire_constant;
    -- logger for split-operator MUX_839_inst flow-through 
    process(IMA82_840) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_839_inst:flowthrough inputs: " & " BITSEL_u8_u1_834_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_834_wire) & " type_cast_836_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_836_wire_constant) & " type_cast_838_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_838_wire_constant) & " outputs:" & " IMA82_840= "  & Convert_SLV_To_Hex_String(IMA82_840));
      --
    end process; 
    -- flow-through select operator MUX_839_inst
    IMA82_840 <= type_cast_836_wire_constant when (BITSEL_u8_u1_834_wire(0) /=  '0') else type_cast_838_wire_constant;
    -- logger for split-operator MUX_849_inst flow-through 
    process(IMA83_850) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_849_inst:flowthrough inputs: " & " BITSEL_u8_u1_844_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_844_wire) & " type_cast_846_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_846_wire_constant) & " type_cast_848_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_848_wire_constant) & " outputs:" & " IMA83_850= "  & Convert_SLV_To_Hex_String(IMA83_850));
      --
    end process; 
    -- flow-through select operator MUX_849_inst
    IMA83_850 <= type_cast_846_wire_constant when (BITSEL_u8_u1_844_wire(0) /=  '0') else type_cast_848_wire_constant;
    -- logger for split-operator MUX_859_inst flow-through 
    process(IMA84_860) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_859_inst:flowthrough inputs: " & " BITSEL_u8_u1_854_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_854_wire) & " type_cast_856_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_856_wire_constant) & " type_cast_858_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_858_wire_constant) & " outputs:" & " IMA84_860= "  & Convert_SLV_To_Hex_String(IMA84_860));
      --
    end process; 
    -- flow-through select operator MUX_859_inst
    IMA84_860 <= type_cast_856_wire_constant when (BITSEL_u8_u1_854_wire(0) /=  '0') else type_cast_858_wire_constant;
    -- logger for split-operator MUX_869_inst flow-through 
    process(IMA85_870) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_869_inst:flowthrough inputs: " & " BITSEL_u8_u1_864_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_864_wire) & " type_cast_866_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_866_wire_constant) & " type_cast_868_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_868_wire_constant) & " outputs:" & " IMA85_870= "  & Convert_SLV_To_Hex_String(IMA85_870));
      --
    end process; 
    -- flow-through select operator MUX_869_inst
    IMA85_870 <= type_cast_866_wire_constant when (BITSEL_u8_u1_864_wire(0) /=  '0') else type_cast_868_wire_constant;
    -- logger for split-operator MUX_879_inst flow-through 
    process(IMA86_880) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_879_inst:flowthrough inputs: " & " BITSEL_u8_u1_874_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_874_wire) & " type_cast_876_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_876_wire_constant) & " type_cast_878_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_878_wire_constant) & " outputs:" & " IMA86_880= "  & Convert_SLV_To_Hex_String(IMA86_880));
      --
    end process; 
    -- flow-through select operator MUX_879_inst
    IMA86_880 <= type_cast_876_wire_constant when (BITSEL_u8_u1_874_wire(0) /=  '0') else type_cast_878_wire_constant;
    -- logger for split-operator MUX_889_inst flow-through 
    process(IMA87_890) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_889_inst:flowthrough inputs: " & " BITSEL_u8_u1_884_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_884_wire) & " type_cast_886_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_886_wire_constant) & " type_cast_888_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_888_wire_constant) & " outputs:" & " IMA87_890= "  & Convert_SLV_To_Hex_String(IMA87_890));
      --
    end process; 
    -- flow-through select operator MUX_889_inst
    IMA87_890 <= type_cast_886_wire_constant when (BITSEL_u8_u1_884_wire(0) /=  '0') else type_cast_888_wire_constant;
    -- logger for split-operator MUX_899_inst flow-through 
    process(IMA88_900) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_899_inst:flowthrough inputs: " & " BITSEL_u8_u1_894_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_894_wire) & " type_cast_896_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_896_wire_constant) & " type_cast_898_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_898_wire_constant) & " outputs:" & " IMA88_900= "  & Convert_SLV_To_Hex_String(IMA88_900));
      --
    end process; 
    -- flow-through select operator MUX_899_inst
    IMA88_900 <= type_cast_896_wire_constant when (BITSEL_u8_u1_894_wire(0) /=  '0') else type_cast_898_wire_constant;
    -- logger for split-operator MUX_89_inst flow-through 
    process(IMA7_90) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_89_inst:flowthrough inputs: " & " BITSEL_u8_u1_84_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_84_wire) & " type_cast_86_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_86_wire_constant) & " type_cast_88_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_88_wire_constant) & " outputs:" & " IMA7_90= "  & Convert_SLV_To_Hex_String(IMA7_90));
      --
    end process; 
    -- flow-through select operator MUX_89_inst
    IMA7_90 <= type_cast_86_wire_constant when (BITSEL_u8_u1_84_wire(0) /=  '0') else type_cast_88_wire_constant;
    -- logger for split-operator MUX_909_inst flow-through 
    process(IMA89_910) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_909_inst:flowthrough inputs: " & " BITSEL_u8_u1_904_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_904_wire) & " type_cast_906_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_906_wire_constant) & " type_cast_908_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_908_wire_constant) & " outputs:" & " IMA89_910= "  & Convert_SLV_To_Hex_String(IMA89_910));
      --
    end process; 
    -- flow-through select operator MUX_909_inst
    IMA89_910 <= type_cast_906_wire_constant when (BITSEL_u8_u1_904_wire(0) /=  '0') else type_cast_908_wire_constant;
    -- logger for split-operator MUX_919_inst flow-through 
    process(IMA90_920) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_919_inst:flowthrough inputs: " & " BITSEL_u8_u1_914_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_914_wire) & " type_cast_916_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_916_wire_constant) & " type_cast_918_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_918_wire_constant) & " outputs:" & " IMA90_920= "  & Convert_SLV_To_Hex_String(IMA90_920));
      --
    end process; 
    -- flow-through select operator MUX_919_inst
    IMA90_920 <= type_cast_916_wire_constant when (BITSEL_u8_u1_914_wire(0) /=  '0') else type_cast_918_wire_constant;
    -- logger for split-operator MUX_929_inst flow-through 
    process(IMA91_930) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_929_inst:flowthrough inputs: " & " BITSEL_u8_u1_924_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_924_wire) & " type_cast_926_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_926_wire_constant) & " type_cast_928_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_928_wire_constant) & " outputs:" & " IMA91_930= "  & Convert_SLV_To_Hex_String(IMA91_930));
      --
    end process; 
    -- flow-through select operator MUX_929_inst
    IMA91_930 <= type_cast_926_wire_constant when (BITSEL_u8_u1_924_wire(0) /=  '0') else type_cast_928_wire_constant;
    -- logger for split-operator MUX_939_inst flow-through 
    process(IMA92_940) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_939_inst:flowthrough inputs: " & " BITSEL_u8_u1_934_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_934_wire) & " type_cast_936_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_936_wire_constant) & " type_cast_938_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_938_wire_constant) & " outputs:" & " IMA92_940= "  & Convert_SLV_To_Hex_String(IMA92_940));
      --
    end process; 
    -- flow-through select operator MUX_939_inst
    IMA92_940 <= type_cast_936_wire_constant when (BITSEL_u8_u1_934_wire(0) /=  '0') else type_cast_938_wire_constant;
    -- logger for split-operator MUX_949_inst flow-through 
    process(IMA93_950) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_949_inst:flowthrough inputs: " & " BITSEL_u8_u1_944_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_944_wire) & " type_cast_946_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_946_wire_constant) & " type_cast_948_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_948_wire_constant) & " outputs:" & " IMA93_950= "  & Convert_SLV_To_Hex_String(IMA93_950));
      --
    end process; 
    -- flow-through select operator MUX_949_inst
    IMA93_950 <= type_cast_946_wire_constant when (BITSEL_u8_u1_944_wire(0) /=  '0') else type_cast_948_wire_constant;
    -- logger for split-operator MUX_959_inst flow-through 
    process(IMA94_960) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_959_inst:flowthrough inputs: " & " BITSEL_u8_u1_954_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_954_wire) & " type_cast_956_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_956_wire_constant) & " type_cast_958_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_958_wire_constant) & " outputs:" & " IMA94_960= "  & Convert_SLV_To_Hex_String(IMA94_960));
      --
    end process; 
    -- flow-through select operator MUX_959_inst
    IMA94_960 <= type_cast_956_wire_constant when (BITSEL_u8_u1_954_wire(0) /=  '0') else type_cast_958_wire_constant;
    -- logger for split-operator MUX_969_inst flow-through 
    process(IMA95_970) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_969_inst:flowthrough inputs: " & " BITSEL_u8_u1_964_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_964_wire) & " type_cast_966_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_966_wire_constant) & " type_cast_968_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_968_wire_constant) & " outputs:" & " IMA95_970= "  & Convert_SLV_To_Hex_String(IMA95_970));
      --
    end process; 
    -- flow-through select operator MUX_969_inst
    IMA95_970 <= type_cast_966_wire_constant when (BITSEL_u8_u1_964_wire(0) /=  '0') else type_cast_968_wire_constant;
    -- logger for split-operator MUX_979_inst flow-through 
    process(IMA96_980) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_979_inst:flowthrough inputs: " & " BITSEL_u8_u1_974_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_974_wire) & " type_cast_976_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_976_wire_constant) & " type_cast_978_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_978_wire_constant) & " outputs:" & " IMA96_980= "  & Convert_SLV_To_Hex_String(IMA96_980));
      --
    end process; 
    -- flow-through select operator MUX_979_inst
    IMA96_980 <= type_cast_976_wire_constant when (BITSEL_u8_u1_974_wire(0) /=  '0') else type_cast_978_wire_constant;
    -- logger for split-operator MUX_989_inst flow-through 
    process(IMA97_990) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_989_inst:flowthrough inputs: " & " BITSEL_u8_u1_984_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_984_wire) & " type_cast_986_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_986_wire_constant) & " type_cast_988_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_988_wire_constant) & " outputs:" & " IMA97_990= "  & Convert_SLV_To_Hex_String(IMA97_990));
      --
    end process; 
    -- flow-through select operator MUX_989_inst
    IMA97_990 <= type_cast_986_wire_constant when (BITSEL_u8_u1_984_wire(0) /=  '0') else type_cast_988_wire_constant;
    -- logger for split-operator MUX_999_inst flow-through 
    process(IMA98_1000) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_999_inst:flowthrough inputs: " & " BITSEL_u8_u1_994_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_994_wire) & " type_cast_996_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_996_wire_constant) & " type_cast_998_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_998_wire_constant) & " outputs:" & " IMA98_1000= "  & Convert_SLV_To_Hex_String(IMA98_1000));
      --
    end process; 
    -- flow-through select operator MUX_999_inst
    IMA98_1000 <= type_cast_996_wire_constant when (BITSEL_u8_u1_994_wire(0) /=  '0') else type_cast_998_wire_constant;
    -- logger for split-operator MUX_99_inst flow-through 
    process(IMA8_100) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:MUX_99_inst:flowthrough inputs: " & " BITSEL_u8_u1_94_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_94_wire) & " type_cast_96_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_96_wire_constant) & " type_cast_98_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_98_wire_constant) & " outputs:" & " IMA8_100= "  & Convert_SLV_To_Hex_String(IMA8_100));
      --
    end process; 
    -- flow-through select operator MUX_99_inst
    IMA8_100 <= type_cast_96_wire_constant when (BITSEL_u8_u1_94_wire(0) /=  '0') else type_cast_98_wire_constant;
    -- logger for split-operator BITSEL_u8_u1_1004_inst flow-through 
    process(BITSEL_u8_u1_1004_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1004_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1003_wire_constant = "& Convert_SLV_To_Hex_String(konst_1003_wire_constant) & " outputs:" & " BITSEL_u8_u1_1004_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1004_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1004_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1003_wire_constant, tmp_var);
      BITSEL_u8_u1_1004_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1014_inst flow-through 
    process(BITSEL_u8_u1_1014_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1014_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1013_wire_constant = "& Convert_SLV_To_Hex_String(konst_1013_wire_constant) & " outputs:" & " BITSEL_u8_u1_1014_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1014_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1014_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1013_wire_constant, tmp_var);
      BITSEL_u8_u1_1014_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1024_inst flow-through 
    process(BITSEL_u8_u1_1024_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1024_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1023_wire_constant = "& Convert_SLV_To_Hex_String(konst_1023_wire_constant) & " outputs:" & " BITSEL_u8_u1_1024_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1024_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1024_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1023_wire_constant, tmp_var);
      BITSEL_u8_u1_1024_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1034_inst flow-through 
    process(BITSEL_u8_u1_1034_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1034_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1033_wire_constant = "& Convert_SLV_To_Hex_String(konst_1033_wire_constant) & " outputs:" & " BITSEL_u8_u1_1034_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1034_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1034_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1033_wire_constant, tmp_var);
      BITSEL_u8_u1_1034_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1044_inst flow-through 
    process(BITSEL_u8_u1_1044_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1044_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1043_wire_constant = "& Convert_SLV_To_Hex_String(konst_1043_wire_constant) & " outputs:" & " BITSEL_u8_u1_1044_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1044_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1044_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1043_wire_constant, tmp_var);
      BITSEL_u8_u1_1044_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_104_inst flow-through 
    process(BITSEL_u8_u1_104_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_104_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_103_wire_constant = "& Convert_SLV_To_Hex_String(konst_103_wire_constant) & " outputs:" & " BITSEL_u8_u1_104_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_104_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_104_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_103_wire_constant, tmp_var);
      BITSEL_u8_u1_104_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1054_inst flow-through 
    process(BITSEL_u8_u1_1054_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1054_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1053_wire_constant = "& Convert_SLV_To_Hex_String(konst_1053_wire_constant) & " outputs:" & " BITSEL_u8_u1_1054_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1054_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1054_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1053_wire_constant, tmp_var);
      BITSEL_u8_u1_1054_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1064_inst flow-through 
    process(BITSEL_u8_u1_1064_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1064_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1063_wire_constant = "& Convert_SLV_To_Hex_String(konst_1063_wire_constant) & " outputs:" & " BITSEL_u8_u1_1064_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1064_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1064_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1063_wire_constant, tmp_var);
      BITSEL_u8_u1_1064_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1074_inst flow-through 
    process(BITSEL_u8_u1_1074_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1074_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1073_wire_constant = "& Convert_SLV_To_Hex_String(konst_1073_wire_constant) & " outputs:" & " BITSEL_u8_u1_1074_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1074_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1074_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1073_wire_constant, tmp_var);
      BITSEL_u8_u1_1074_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1084_inst flow-through 
    process(BITSEL_u8_u1_1084_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1084_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1083_wire_constant = "& Convert_SLV_To_Hex_String(konst_1083_wire_constant) & " outputs:" & " BITSEL_u8_u1_1084_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1084_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1084_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1083_wire_constant, tmp_var);
      BITSEL_u8_u1_1084_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1094_inst flow-through 
    process(BITSEL_u8_u1_1094_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1094_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1093_wire_constant = "& Convert_SLV_To_Hex_String(konst_1093_wire_constant) & " outputs:" & " BITSEL_u8_u1_1094_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1094_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1094_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1093_wire_constant, tmp_var);
      BITSEL_u8_u1_1094_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1104_inst flow-through 
    process(BITSEL_u8_u1_1104_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1104_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1103_wire_constant = "& Convert_SLV_To_Hex_String(konst_1103_wire_constant) & " outputs:" & " BITSEL_u8_u1_1104_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1104_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1104_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1103_wire_constant, tmp_var);
      BITSEL_u8_u1_1104_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1114_inst flow-through 
    process(BITSEL_u8_u1_1114_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1114_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1113_wire_constant = "& Convert_SLV_To_Hex_String(konst_1113_wire_constant) & " outputs:" & " BITSEL_u8_u1_1114_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1114_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1114_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1113_wire_constant, tmp_var);
      BITSEL_u8_u1_1114_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1124_inst flow-through 
    process(BITSEL_u8_u1_1124_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1124_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1123_wire_constant = "& Convert_SLV_To_Hex_String(konst_1123_wire_constant) & " outputs:" & " BITSEL_u8_u1_1124_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1124_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1124_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1123_wire_constant, tmp_var);
      BITSEL_u8_u1_1124_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1134_inst flow-through 
    process(BITSEL_u8_u1_1134_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1134_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1133_wire_constant = "& Convert_SLV_To_Hex_String(konst_1133_wire_constant) & " outputs:" & " BITSEL_u8_u1_1134_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1134_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1134_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1133_wire_constant, tmp_var);
      BITSEL_u8_u1_1134_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1144_inst flow-through 
    process(BITSEL_u8_u1_1144_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1144_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1143_wire_constant = "& Convert_SLV_To_Hex_String(konst_1143_wire_constant) & " outputs:" & " BITSEL_u8_u1_1144_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1144_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1144_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1143_wire_constant, tmp_var);
      BITSEL_u8_u1_1144_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_114_inst flow-through 
    process(BITSEL_u8_u1_114_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_114_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_113_wire_constant = "& Convert_SLV_To_Hex_String(konst_113_wire_constant) & " outputs:" & " BITSEL_u8_u1_114_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_114_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_114_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_113_wire_constant, tmp_var);
      BITSEL_u8_u1_114_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1154_inst flow-through 
    process(BITSEL_u8_u1_1154_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1154_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1153_wire_constant = "& Convert_SLV_To_Hex_String(konst_1153_wire_constant) & " outputs:" & " BITSEL_u8_u1_1154_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1154_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1154_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1153_wire_constant, tmp_var);
      BITSEL_u8_u1_1154_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1164_inst flow-through 
    process(BITSEL_u8_u1_1164_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1164_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1163_wire_constant = "& Convert_SLV_To_Hex_String(konst_1163_wire_constant) & " outputs:" & " BITSEL_u8_u1_1164_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1164_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1164_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1163_wire_constant, tmp_var);
      BITSEL_u8_u1_1164_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1174_inst flow-through 
    process(BITSEL_u8_u1_1174_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1174_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1173_wire_constant = "& Convert_SLV_To_Hex_String(konst_1173_wire_constant) & " outputs:" & " BITSEL_u8_u1_1174_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1174_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1174_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1173_wire_constant, tmp_var);
      BITSEL_u8_u1_1174_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1184_inst flow-through 
    process(BITSEL_u8_u1_1184_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1184_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1183_wire_constant = "& Convert_SLV_To_Hex_String(konst_1183_wire_constant) & " outputs:" & " BITSEL_u8_u1_1184_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1184_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1184_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1183_wire_constant, tmp_var);
      BITSEL_u8_u1_1184_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1194_inst flow-through 
    process(BITSEL_u8_u1_1194_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1194_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1193_wire_constant = "& Convert_SLV_To_Hex_String(konst_1193_wire_constant) & " outputs:" & " BITSEL_u8_u1_1194_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1194_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1194_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1193_wire_constant, tmp_var);
      BITSEL_u8_u1_1194_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1204_inst flow-through 
    process(BITSEL_u8_u1_1204_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1204_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1203_wire_constant = "& Convert_SLV_To_Hex_String(konst_1203_wire_constant) & " outputs:" & " BITSEL_u8_u1_1204_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1204_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1204_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1203_wire_constant, tmp_var);
      BITSEL_u8_u1_1204_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1214_inst flow-through 
    process(BITSEL_u8_u1_1214_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1214_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1213_wire_constant = "& Convert_SLV_To_Hex_String(konst_1213_wire_constant) & " outputs:" & " BITSEL_u8_u1_1214_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1214_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1214_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1213_wire_constant, tmp_var);
      BITSEL_u8_u1_1214_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1224_inst flow-through 
    process(BITSEL_u8_u1_1224_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1224_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1223_wire_constant = "& Convert_SLV_To_Hex_String(konst_1223_wire_constant) & " outputs:" & " BITSEL_u8_u1_1224_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1224_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1224_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1223_wire_constant, tmp_var);
      BITSEL_u8_u1_1224_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1234_inst flow-through 
    process(BITSEL_u8_u1_1234_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1234_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1233_wire_constant = "& Convert_SLV_To_Hex_String(konst_1233_wire_constant) & " outputs:" & " BITSEL_u8_u1_1234_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1234_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1234_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1233_wire_constant, tmp_var);
      BITSEL_u8_u1_1234_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1244_inst flow-through 
    process(BITSEL_u8_u1_1244_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1244_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1243_wire_constant = "& Convert_SLV_To_Hex_String(konst_1243_wire_constant) & " outputs:" & " BITSEL_u8_u1_1244_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1244_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1244_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1243_wire_constant, tmp_var);
      BITSEL_u8_u1_1244_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_124_inst flow-through 
    process(BITSEL_u8_u1_124_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_124_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_123_wire_constant = "& Convert_SLV_To_Hex_String(konst_123_wire_constant) & " outputs:" & " BITSEL_u8_u1_124_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_124_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_124_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_123_wire_constant, tmp_var);
      BITSEL_u8_u1_124_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1254_inst flow-through 
    process(BITSEL_u8_u1_1254_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1254_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1253_wire_constant = "& Convert_SLV_To_Hex_String(konst_1253_wire_constant) & " outputs:" & " BITSEL_u8_u1_1254_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1254_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1254_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1253_wire_constant, tmp_var);
      BITSEL_u8_u1_1254_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1264_inst flow-through 
    process(BITSEL_u8_u1_1264_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1264_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1263_wire_constant = "& Convert_SLV_To_Hex_String(konst_1263_wire_constant) & " outputs:" & " BITSEL_u8_u1_1264_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1264_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1264_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1263_wire_constant, tmp_var);
      BITSEL_u8_u1_1264_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1274_inst flow-through 
    process(BITSEL_u8_u1_1274_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1274_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1273_wire_constant = "& Convert_SLV_To_Hex_String(konst_1273_wire_constant) & " outputs:" & " BITSEL_u8_u1_1274_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1274_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1274_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1273_wire_constant, tmp_var);
      BITSEL_u8_u1_1274_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1284_inst flow-through 
    process(BITSEL_u8_u1_1284_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1284_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1283_wire_constant = "& Convert_SLV_To_Hex_String(konst_1283_wire_constant) & " outputs:" & " BITSEL_u8_u1_1284_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1284_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1284_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1283_wire_constant, tmp_var);
      BITSEL_u8_u1_1284_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1294_inst flow-through 
    process(BITSEL_u8_u1_1294_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1294_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1293_wire_constant = "& Convert_SLV_To_Hex_String(konst_1293_wire_constant) & " outputs:" & " BITSEL_u8_u1_1294_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1294_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1294_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1293_wire_constant, tmp_var);
      BITSEL_u8_u1_1294_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1302_inst flow-through 
    process(BITSEL_u8_u1_1302_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1302_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1301_wire_constant = "& Convert_SLV_To_Hex_String(konst_1301_wire_constant) & " outputs:" & " BITSEL_u8_u1_1302_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1302_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1302_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1301_wire_constant, tmp_var);
      BITSEL_u8_u1_1302_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1310_inst flow-through 
    process(BITSEL_u8_u1_1310_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1310_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1309_wire_constant = "& Convert_SLV_To_Hex_String(konst_1309_wire_constant) & " outputs:" & " BITSEL_u8_u1_1310_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1310_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1310_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1309_wire_constant, tmp_var);
      BITSEL_u8_u1_1310_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1318_inst flow-through 
    process(BITSEL_u8_u1_1318_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1318_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1317_wire_constant = "& Convert_SLV_To_Hex_String(konst_1317_wire_constant) & " outputs:" & " BITSEL_u8_u1_1318_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1318_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1318_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1317_wire_constant, tmp_var);
      BITSEL_u8_u1_1318_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1326_inst flow-through 
    process(BITSEL_u8_u1_1326_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1326_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1325_wire_constant = "& Convert_SLV_To_Hex_String(konst_1325_wire_constant) & " outputs:" & " BITSEL_u8_u1_1326_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1326_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1326_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1325_wire_constant, tmp_var);
      BITSEL_u8_u1_1326_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1334_inst flow-through 
    process(BITSEL_u8_u1_1334_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1334_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1333_wire_constant = "& Convert_SLV_To_Hex_String(konst_1333_wire_constant) & " outputs:" & " BITSEL_u8_u1_1334_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1334_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1334_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1333_wire_constant, tmp_var);
      BITSEL_u8_u1_1334_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1342_inst flow-through 
    process(BITSEL_u8_u1_1342_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1342_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1341_wire_constant = "& Convert_SLV_To_Hex_String(konst_1341_wire_constant) & " outputs:" & " BITSEL_u8_u1_1342_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1342_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1342_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1341_wire_constant, tmp_var);
      BITSEL_u8_u1_1342_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_134_inst flow-through 
    process(BITSEL_u8_u1_134_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_134_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_133_wire_constant = "& Convert_SLV_To_Hex_String(konst_133_wire_constant) & " outputs:" & " BITSEL_u8_u1_134_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_134_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_134_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_133_wire_constant, tmp_var);
      BITSEL_u8_u1_134_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1350_inst flow-through 
    process(BITSEL_u8_u1_1350_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1350_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1349_wire_constant = "& Convert_SLV_To_Hex_String(konst_1349_wire_constant) & " outputs:" & " BITSEL_u8_u1_1350_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1350_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1350_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1349_wire_constant, tmp_var);
      BITSEL_u8_u1_1350_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1358_inst flow-through 
    process(BITSEL_u8_u1_1358_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1358_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1357_wire_constant = "& Convert_SLV_To_Hex_String(konst_1357_wire_constant) & " outputs:" & " BITSEL_u8_u1_1358_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1358_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1358_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1357_wire_constant, tmp_var);
      BITSEL_u8_u1_1358_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1366_inst flow-through 
    process(BITSEL_u8_u1_1366_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1366_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1365_wire_constant = "& Convert_SLV_To_Hex_String(konst_1365_wire_constant) & " outputs:" & " BITSEL_u8_u1_1366_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1366_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1366_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1365_wire_constant, tmp_var);
      BITSEL_u8_u1_1366_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1374_inst flow-through 
    process(BITSEL_u8_u1_1374_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1374_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1373_wire_constant = "& Convert_SLV_To_Hex_String(konst_1373_wire_constant) & " outputs:" & " BITSEL_u8_u1_1374_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1374_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1374_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1373_wire_constant, tmp_var);
      BITSEL_u8_u1_1374_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1382_inst flow-through 
    process(BITSEL_u8_u1_1382_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1382_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1381_wire_constant = "& Convert_SLV_To_Hex_String(konst_1381_wire_constant) & " outputs:" & " BITSEL_u8_u1_1382_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1382_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1382_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1381_wire_constant, tmp_var);
      BITSEL_u8_u1_1382_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1390_inst flow-through 
    process(BITSEL_u8_u1_1390_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1390_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1389_wire_constant = "& Convert_SLV_To_Hex_String(konst_1389_wire_constant) & " outputs:" & " BITSEL_u8_u1_1390_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1390_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1390_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1389_wire_constant, tmp_var);
      BITSEL_u8_u1_1390_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1398_inst flow-through 
    process(BITSEL_u8_u1_1398_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1398_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1397_wire_constant = "& Convert_SLV_To_Hex_String(konst_1397_wire_constant) & " outputs:" & " BITSEL_u8_u1_1398_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1398_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1398_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1397_wire_constant, tmp_var);
      BITSEL_u8_u1_1398_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_13_inst flow-through 
    process(BITSEL_u8_u1_13_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_13_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_12_wire_constant = "& Convert_SLV_To_Hex_String(konst_12_wire_constant) & " outputs:" & " BITSEL_u8_u1_13_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_13_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_13_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_12_wire_constant, tmp_var);
      BITSEL_u8_u1_13_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1406_inst flow-through 
    process(BITSEL_u8_u1_1406_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1406_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1405_wire_constant = "& Convert_SLV_To_Hex_String(konst_1405_wire_constant) & " outputs:" & " BITSEL_u8_u1_1406_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1406_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1406_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1405_wire_constant, tmp_var);
      BITSEL_u8_u1_1406_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1414_inst flow-through 
    process(BITSEL_u8_u1_1414_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1414_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1413_wire_constant = "& Convert_SLV_To_Hex_String(konst_1413_wire_constant) & " outputs:" & " BITSEL_u8_u1_1414_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1414_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1414_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1413_wire_constant, tmp_var);
      BITSEL_u8_u1_1414_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1422_inst flow-through 
    process(BITSEL_u8_u1_1422_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1422_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1421_wire_constant = "& Convert_SLV_To_Hex_String(konst_1421_wire_constant) & " outputs:" & " BITSEL_u8_u1_1422_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1422_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1422_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1421_wire_constant, tmp_var);
      BITSEL_u8_u1_1422_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1430_inst flow-through 
    process(BITSEL_u8_u1_1430_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1430_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1429_wire_constant = "& Convert_SLV_To_Hex_String(konst_1429_wire_constant) & " outputs:" & " BITSEL_u8_u1_1430_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1430_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1430_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1429_wire_constant, tmp_var);
      BITSEL_u8_u1_1430_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1438_inst flow-through 
    process(BITSEL_u8_u1_1438_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1438_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1437_wire_constant = "& Convert_SLV_To_Hex_String(konst_1437_wire_constant) & " outputs:" & " BITSEL_u8_u1_1438_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1438_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1438_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1437_wire_constant, tmp_var);
      BITSEL_u8_u1_1438_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1446_inst flow-through 
    process(BITSEL_u8_u1_1446_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1446_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1445_wire_constant = "& Convert_SLV_To_Hex_String(konst_1445_wire_constant) & " outputs:" & " BITSEL_u8_u1_1446_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1446_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1446_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1445_wire_constant, tmp_var);
      BITSEL_u8_u1_1446_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_144_inst flow-through 
    process(BITSEL_u8_u1_144_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_144_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_143_wire_constant = "& Convert_SLV_To_Hex_String(konst_143_wire_constant) & " outputs:" & " BITSEL_u8_u1_144_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_144_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_144_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_143_wire_constant, tmp_var);
      BITSEL_u8_u1_144_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1454_inst flow-through 
    process(BITSEL_u8_u1_1454_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1454_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1453_wire_constant = "& Convert_SLV_To_Hex_String(konst_1453_wire_constant) & " outputs:" & " BITSEL_u8_u1_1454_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1454_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1454_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1453_wire_constant, tmp_var);
      BITSEL_u8_u1_1454_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1462_inst flow-through 
    process(BITSEL_u8_u1_1462_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1462_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1461_wire_constant = "& Convert_SLV_To_Hex_String(konst_1461_wire_constant) & " outputs:" & " BITSEL_u8_u1_1462_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1462_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1462_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1461_wire_constant, tmp_var);
      BITSEL_u8_u1_1462_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1470_inst flow-through 
    process(BITSEL_u8_u1_1470_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1470_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1469_wire_constant = "& Convert_SLV_To_Hex_String(konst_1469_wire_constant) & " outputs:" & " BITSEL_u8_u1_1470_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1470_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1470_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1469_wire_constant, tmp_var);
      BITSEL_u8_u1_1470_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1478_inst flow-through 
    process(BITSEL_u8_u1_1478_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1478_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1477_wire_constant = "& Convert_SLV_To_Hex_String(konst_1477_wire_constant) & " outputs:" & " BITSEL_u8_u1_1478_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1478_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1478_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1477_wire_constant, tmp_var);
      BITSEL_u8_u1_1478_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1486_inst flow-through 
    process(BITSEL_u8_u1_1486_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1486_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1485_wire_constant = "& Convert_SLV_To_Hex_String(konst_1485_wire_constant) & " outputs:" & " BITSEL_u8_u1_1486_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1486_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1486_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1485_wire_constant, tmp_var);
      BITSEL_u8_u1_1486_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1494_inst flow-through 
    process(BITSEL_u8_u1_1494_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1494_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1493_wire_constant = "& Convert_SLV_To_Hex_String(konst_1493_wire_constant) & " outputs:" & " BITSEL_u8_u1_1494_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1494_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1494_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1493_wire_constant, tmp_var);
      BITSEL_u8_u1_1494_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1502_inst flow-through 
    process(BITSEL_u8_u1_1502_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1502_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1501_wire_constant = "& Convert_SLV_To_Hex_String(konst_1501_wire_constant) & " outputs:" & " BITSEL_u8_u1_1502_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1502_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1502_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1501_wire_constant, tmp_var);
      BITSEL_u8_u1_1502_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1510_inst flow-through 
    process(BITSEL_u8_u1_1510_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1510_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1509_wire_constant = "& Convert_SLV_To_Hex_String(konst_1509_wire_constant) & " outputs:" & " BITSEL_u8_u1_1510_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1510_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1510_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1509_wire_constant, tmp_var);
      BITSEL_u8_u1_1510_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1518_inst flow-through 
    process(BITSEL_u8_u1_1518_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1518_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1517_wire_constant = "& Convert_SLV_To_Hex_String(konst_1517_wire_constant) & " outputs:" & " BITSEL_u8_u1_1518_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1518_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1518_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1517_wire_constant, tmp_var);
      BITSEL_u8_u1_1518_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1526_inst flow-through 
    process(BITSEL_u8_u1_1526_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1526_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1525_wire_constant = "& Convert_SLV_To_Hex_String(konst_1525_wire_constant) & " outputs:" & " BITSEL_u8_u1_1526_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1526_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1526_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1525_wire_constant, tmp_var);
      BITSEL_u8_u1_1526_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1534_inst flow-through 
    process(BITSEL_u8_u1_1534_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1534_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1533_wire_constant = "& Convert_SLV_To_Hex_String(konst_1533_wire_constant) & " outputs:" & " BITSEL_u8_u1_1534_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1534_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1534_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1533_wire_constant, tmp_var);
      BITSEL_u8_u1_1534_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1542_inst flow-through 
    process(BITSEL_u8_u1_1542_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1542_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1541_wire_constant = "& Convert_SLV_To_Hex_String(konst_1541_wire_constant) & " outputs:" & " BITSEL_u8_u1_1542_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1542_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1542_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1541_wire_constant, tmp_var);
      BITSEL_u8_u1_1542_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_154_inst flow-through 
    process(BITSEL_u8_u1_154_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_154_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_153_wire_constant = "& Convert_SLV_To_Hex_String(konst_153_wire_constant) & " outputs:" & " BITSEL_u8_u1_154_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_154_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_154_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_153_wire_constant, tmp_var);
      BITSEL_u8_u1_154_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1550_inst flow-through 
    process(BITSEL_u8_u1_1550_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1550_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1549_wire_constant = "& Convert_SLV_To_Hex_String(konst_1549_wire_constant) & " outputs:" & " BITSEL_u8_u1_1550_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1550_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1550_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1549_wire_constant, tmp_var);
      BITSEL_u8_u1_1550_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1558_inst flow-through 
    process(BITSEL_u8_u1_1558_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1558_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1557_wire_constant = "& Convert_SLV_To_Hex_String(konst_1557_wire_constant) & " outputs:" & " BITSEL_u8_u1_1558_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1558_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1558_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1557_wire_constant, tmp_var);
      BITSEL_u8_u1_1558_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1566_inst flow-through 
    process(BITSEL_u8_u1_1566_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1566_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1565_wire_constant = "& Convert_SLV_To_Hex_String(konst_1565_wire_constant) & " outputs:" & " BITSEL_u8_u1_1566_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1566_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1566_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1565_wire_constant, tmp_var);
      BITSEL_u8_u1_1566_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1574_inst flow-through 
    process(BITSEL_u8_u1_1574_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1574_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1573_wire_constant = "& Convert_SLV_To_Hex_String(konst_1573_wire_constant) & " outputs:" & " BITSEL_u8_u1_1574_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1574_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1574_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1573_wire_constant, tmp_var);
      BITSEL_u8_u1_1574_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1582_inst flow-through 
    process(BITSEL_u8_u1_1582_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1582_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1581_wire_constant = "& Convert_SLV_To_Hex_String(konst_1581_wire_constant) & " outputs:" & " BITSEL_u8_u1_1582_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1582_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1582_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1581_wire_constant, tmp_var);
      BITSEL_u8_u1_1582_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1590_inst flow-through 
    process(BITSEL_u8_u1_1590_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1590_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1589_wire_constant = "& Convert_SLV_To_Hex_String(konst_1589_wire_constant) & " outputs:" & " BITSEL_u8_u1_1590_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1590_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1590_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1589_wire_constant, tmp_var);
      BITSEL_u8_u1_1590_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1598_inst flow-through 
    process(BITSEL_u8_u1_1598_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1598_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1597_wire_constant = "& Convert_SLV_To_Hex_String(konst_1597_wire_constant) & " outputs:" & " BITSEL_u8_u1_1598_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1598_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1598_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1597_wire_constant, tmp_var);
      BITSEL_u8_u1_1598_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1606_inst flow-through 
    process(BITSEL_u8_u1_1606_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1606_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1605_wire_constant = "& Convert_SLV_To_Hex_String(konst_1605_wire_constant) & " outputs:" & " BITSEL_u8_u1_1606_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1606_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1606_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1605_wire_constant, tmp_var);
      BITSEL_u8_u1_1606_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1614_inst flow-through 
    process(BITSEL_u8_u1_1614_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1614_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1613_wire_constant = "& Convert_SLV_To_Hex_String(konst_1613_wire_constant) & " outputs:" & " BITSEL_u8_u1_1614_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1614_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1614_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1613_wire_constant, tmp_var);
      BITSEL_u8_u1_1614_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1622_inst flow-through 
    process(BITSEL_u8_u1_1622_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1622_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1621_wire_constant = "& Convert_SLV_To_Hex_String(konst_1621_wire_constant) & " outputs:" & " BITSEL_u8_u1_1622_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1622_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1622_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1621_wire_constant, tmp_var);
      BITSEL_u8_u1_1622_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1630_inst flow-through 
    process(BITSEL_u8_u1_1630_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1630_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1629_wire_constant = "& Convert_SLV_To_Hex_String(konst_1629_wire_constant) & " outputs:" & " BITSEL_u8_u1_1630_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1630_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1630_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1629_wire_constant, tmp_var);
      BITSEL_u8_u1_1630_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1638_inst flow-through 
    process(BITSEL_u8_u1_1638_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1638_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1637_wire_constant = "& Convert_SLV_To_Hex_String(konst_1637_wire_constant) & " outputs:" & " BITSEL_u8_u1_1638_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1638_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1638_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1637_wire_constant, tmp_var);
      BITSEL_u8_u1_1638_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1646_inst flow-through 
    process(BITSEL_u8_u1_1646_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1646_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1645_wire_constant = "& Convert_SLV_To_Hex_String(konst_1645_wire_constant) & " outputs:" & " BITSEL_u8_u1_1646_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1646_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1646_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1645_wire_constant, tmp_var);
      BITSEL_u8_u1_1646_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_164_inst flow-through 
    process(BITSEL_u8_u1_164_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_164_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_163_wire_constant = "& Convert_SLV_To_Hex_String(konst_163_wire_constant) & " outputs:" & " BITSEL_u8_u1_164_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_164_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_164_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_163_wire_constant, tmp_var);
      BITSEL_u8_u1_164_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1654_inst flow-through 
    process(BITSEL_u8_u1_1654_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1654_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1653_wire_constant = "& Convert_SLV_To_Hex_String(konst_1653_wire_constant) & " outputs:" & " BITSEL_u8_u1_1654_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1654_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1654_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1653_wire_constant, tmp_var);
      BITSEL_u8_u1_1654_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1662_inst flow-through 
    process(BITSEL_u8_u1_1662_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1662_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1661_wire_constant = "& Convert_SLV_To_Hex_String(konst_1661_wire_constant) & " outputs:" & " BITSEL_u8_u1_1662_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1662_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1662_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1661_wire_constant, tmp_var);
      BITSEL_u8_u1_1662_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1670_inst flow-through 
    process(BITSEL_u8_u1_1670_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1670_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1669_wire_constant = "& Convert_SLV_To_Hex_String(konst_1669_wire_constant) & " outputs:" & " BITSEL_u8_u1_1670_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1670_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1670_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1669_wire_constant, tmp_var);
      BITSEL_u8_u1_1670_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1678_inst flow-through 
    process(BITSEL_u8_u1_1678_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1678_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1677_wire_constant = "& Convert_SLV_To_Hex_String(konst_1677_wire_constant) & " outputs:" & " BITSEL_u8_u1_1678_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1678_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1678_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1677_wire_constant, tmp_var);
      BITSEL_u8_u1_1678_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1686_inst flow-through 
    process(BITSEL_u8_u1_1686_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1686_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1685_wire_constant = "& Convert_SLV_To_Hex_String(konst_1685_wire_constant) & " outputs:" & " BITSEL_u8_u1_1686_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1686_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1686_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1685_wire_constant, tmp_var);
      BITSEL_u8_u1_1686_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1694_inst flow-through 
    process(BITSEL_u8_u1_1694_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1694_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1693_wire_constant = "& Convert_SLV_To_Hex_String(konst_1693_wire_constant) & " outputs:" & " BITSEL_u8_u1_1694_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1694_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1694_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1693_wire_constant, tmp_var);
      BITSEL_u8_u1_1694_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1702_inst flow-through 
    process(BITSEL_u8_u1_1702_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1702_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1701_wire_constant = "& Convert_SLV_To_Hex_String(konst_1701_wire_constant) & " outputs:" & " BITSEL_u8_u1_1702_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1702_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1702_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1701_wire_constant, tmp_var);
      BITSEL_u8_u1_1702_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1710_inst flow-through 
    process(BITSEL_u8_u1_1710_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1710_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1709_wire_constant = "& Convert_SLV_To_Hex_String(konst_1709_wire_constant) & " outputs:" & " BITSEL_u8_u1_1710_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1710_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1710_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1709_wire_constant, tmp_var);
      BITSEL_u8_u1_1710_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1718_inst flow-through 
    process(BITSEL_u8_u1_1718_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1718_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1717_wire_constant = "& Convert_SLV_To_Hex_String(konst_1717_wire_constant) & " outputs:" & " BITSEL_u8_u1_1718_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1718_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1718_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1717_wire_constant, tmp_var);
      BITSEL_u8_u1_1718_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1726_inst flow-through 
    process(BITSEL_u8_u1_1726_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1726_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1725_wire_constant = "& Convert_SLV_To_Hex_String(konst_1725_wire_constant) & " outputs:" & " BITSEL_u8_u1_1726_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1726_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1726_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1725_wire_constant, tmp_var);
      BITSEL_u8_u1_1726_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1734_inst flow-through 
    process(BITSEL_u8_u1_1734_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1734_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1733_wire_constant = "& Convert_SLV_To_Hex_String(konst_1733_wire_constant) & " outputs:" & " BITSEL_u8_u1_1734_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1734_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1734_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1733_wire_constant, tmp_var);
      BITSEL_u8_u1_1734_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1742_inst flow-through 
    process(BITSEL_u8_u1_1742_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1742_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1741_wire_constant = "& Convert_SLV_To_Hex_String(konst_1741_wire_constant) & " outputs:" & " BITSEL_u8_u1_1742_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1742_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1742_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1741_wire_constant, tmp_var);
      BITSEL_u8_u1_1742_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_174_inst flow-through 
    process(BITSEL_u8_u1_174_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_174_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_173_wire_constant = "& Convert_SLV_To_Hex_String(konst_173_wire_constant) & " outputs:" & " BITSEL_u8_u1_174_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_174_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_174_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_173_wire_constant, tmp_var);
      BITSEL_u8_u1_174_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1750_inst flow-through 
    process(BITSEL_u8_u1_1750_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1750_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1749_wire_constant = "& Convert_SLV_To_Hex_String(konst_1749_wire_constant) & " outputs:" & " BITSEL_u8_u1_1750_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1750_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1750_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1749_wire_constant, tmp_var);
      BITSEL_u8_u1_1750_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1758_inst flow-through 
    process(BITSEL_u8_u1_1758_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1758_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1757_wire_constant = "& Convert_SLV_To_Hex_String(konst_1757_wire_constant) & " outputs:" & " BITSEL_u8_u1_1758_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1758_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1758_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1757_wire_constant, tmp_var);
      BITSEL_u8_u1_1758_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1766_inst flow-through 
    process(BITSEL_u8_u1_1766_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1766_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1765_wire_constant = "& Convert_SLV_To_Hex_String(konst_1765_wire_constant) & " outputs:" & " BITSEL_u8_u1_1766_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1766_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1766_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1765_wire_constant, tmp_var);
      BITSEL_u8_u1_1766_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1774_inst flow-through 
    process(BITSEL_u8_u1_1774_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1774_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1773_wire_constant = "& Convert_SLV_To_Hex_String(konst_1773_wire_constant) & " outputs:" & " BITSEL_u8_u1_1774_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1774_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1774_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1773_wire_constant, tmp_var);
      BITSEL_u8_u1_1774_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1782_inst flow-through 
    process(BITSEL_u8_u1_1782_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1782_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1781_wire_constant = "& Convert_SLV_To_Hex_String(konst_1781_wire_constant) & " outputs:" & " BITSEL_u8_u1_1782_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1782_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1782_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1781_wire_constant, tmp_var);
      BITSEL_u8_u1_1782_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1790_inst flow-through 
    process(BITSEL_u8_u1_1790_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1790_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1789_wire_constant = "& Convert_SLV_To_Hex_String(konst_1789_wire_constant) & " outputs:" & " BITSEL_u8_u1_1790_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1790_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1790_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1789_wire_constant, tmp_var);
      BITSEL_u8_u1_1790_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1798_inst flow-through 
    process(BITSEL_u8_u1_1798_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1798_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1797_wire_constant = "& Convert_SLV_To_Hex_String(konst_1797_wire_constant) & " outputs:" & " BITSEL_u8_u1_1798_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1798_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1798_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1797_wire_constant, tmp_var);
      BITSEL_u8_u1_1798_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1806_inst flow-through 
    process(BITSEL_u8_u1_1806_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1806_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1805_wire_constant = "& Convert_SLV_To_Hex_String(konst_1805_wire_constant) & " outputs:" & " BITSEL_u8_u1_1806_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1806_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1806_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1805_wire_constant, tmp_var);
      BITSEL_u8_u1_1806_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1814_inst flow-through 
    process(BITSEL_u8_u1_1814_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1814_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1813_wire_constant = "& Convert_SLV_To_Hex_String(konst_1813_wire_constant) & " outputs:" & " BITSEL_u8_u1_1814_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1814_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1814_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1813_wire_constant, tmp_var);
      BITSEL_u8_u1_1814_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1822_inst flow-through 
    process(BITSEL_u8_u1_1822_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1822_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1821_wire_constant = "& Convert_SLV_To_Hex_String(konst_1821_wire_constant) & " outputs:" & " BITSEL_u8_u1_1822_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1822_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1822_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1821_wire_constant, tmp_var);
      BITSEL_u8_u1_1822_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1830_inst flow-through 
    process(BITSEL_u8_u1_1830_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1830_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1829_wire_constant = "& Convert_SLV_To_Hex_String(konst_1829_wire_constant) & " outputs:" & " BITSEL_u8_u1_1830_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1830_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1830_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1829_wire_constant, tmp_var);
      BITSEL_u8_u1_1830_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1838_inst flow-through 
    process(BITSEL_u8_u1_1838_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1838_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1837_wire_constant = "& Convert_SLV_To_Hex_String(konst_1837_wire_constant) & " outputs:" & " BITSEL_u8_u1_1838_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1838_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1838_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1837_wire_constant, tmp_var);
      BITSEL_u8_u1_1838_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1846_inst flow-through 
    process(BITSEL_u8_u1_1846_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1846_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1845_wire_constant = "& Convert_SLV_To_Hex_String(konst_1845_wire_constant) & " outputs:" & " BITSEL_u8_u1_1846_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1846_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1846_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1845_wire_constant, tmp_var);
      BITSEL_u8_u1_1846_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_184_inst flow-through 
    process(BITSEL_u8_u1_184_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_184_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_183_wire_constant = "& Convert_SLV_To_Hex_String(konst_183_wire_constant) & " outputs:" & " BITSEL_u8_u1_184_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_184_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_184_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_183_wire_constant, tmp_var);
      BITSEL_u8_u1_184_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1854_inst flow-through 
    process(BITSEL_u8_u1_1854_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1854_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1853_wire_constant = "& Convert_SLV_To_Hex_String(konst_1853_wire_constant) & " outputs:" & " BITSEL_u8_u1_1854_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1854_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1854_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1853_wire_constant, tmp_var);
      BITSEL_u8_u1_1854_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1862_inst flow-through 
    process(BITSEL_u8_u1_1862_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1862_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1861_wire_constant = "& Convert_SLV_To_Hex_String(konst_1861_wire_constant) & " outputs:" & " BITSEL_u8_u1_1862_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1862_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1862_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1861_wire_constant, tmp_var);
      BITSEL_u8_u1_1862_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1870_inst flow-through 
    process(BITSEL_u8_u1_1870_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1870_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1869_wire_constant = "& Convert_SLV_To_Hex_String(konst_1869_wire_constant) & " outputs:" & " BITSEL_u8_u1_1870_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1870_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1870_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1869_wire_constant, tmp_var);
      BITSEL_u8_u1_1870_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1878_inst flow-through 
    process(BITSEL_u8_u1_1878_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1878_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1877_wire_constant = "& Convert_SLV_To_Hex_String(konst_1877_wire_constant) & " outputs:" & " BITSEL_u8_u1_1878_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1878_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1878_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1877_wire_constant, tmp_var);
      BITSEL_u8_u1_1878_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1886_inst flow-through 
    process(BITSEL_u8_u1_1886_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1886_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1885_wire_constant = "& Convert_SLV_To_Hex_String(konst_1885_wire_constant) & " outputs:" & " BITSEL_u8_u1_1886_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1886_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1886_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1885_wire_constant, tmp_var);
      BITSEL_u8_u1_1886_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1894_inst flow-through 
    process(BITSEL_u8_u1_1894_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1894_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1893_wire_constant = "& Convert_SLV_To_Hex_String(konst_1893_wire_constant) & " outputs:" & " BITSEL_u8_u1_1894_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1894_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1894_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1893_wire_constant, tmp_var);
      BITSEL_u8_u1_1894_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1902_inst flow-through 
    process(BITSEL_u8_u1_1902_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1902_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1901_wire_constant = "& Convert_SLV_To_Hex_String(konst_1901_wire_constant) & " outputs:" & " BITSEL_u8_u1_1902_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1902_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1902_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1901_wire_constant, tmp_var);
      BITSEL_u8_u1_1902_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1910_inst flow-through 
    process(BITSEL_u8_u1_1910_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1910_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1909_wire_constant = "& Convert_SLV_To_Hex_String(konst_1909_wire_constant) & " outputs:" & " BITSEL_u8_u1_1910_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1910_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1910_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1909_wire_constant, tmp_var);
      BITSEL_u8_u1_1910_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1918_inst flow-through 
    process(BITSEL_u8_u1_1918_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1918_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1917_wire_constant = "& Convert_SLV_To_Hex_String(konst_1917_wire_constant) & " outputs:" & " BITSEL_u8_u1_1918_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1918_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1918_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1917_wire_constant, tmp_var);
      BITSEL_u8_u1_1918_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1926_inst flow-through 
    process(BITSEL_u8_u1_1926_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1926_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1925_wire_constant = "& Convert_SLV_To_Hex_String(konst_1925_wire_constant) & " outputs:" & " BITSEL_u8_u1_1926_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1926_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1926_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1925_wire_constant, tmp_var);
      BITSEL_u8_u1_1926_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1934_inst flow-through 
    process(BITSEL_u8_u1_1934_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1934_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1933_wire_constant = "& Convert_SLV_To_Hex_String(konst_1933_wire_constant) & " outputs:" & " BITSEL_u8_u1_1934_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1934_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1934_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1933_wire_constant, tmp_var);
      BITSEL_u8_u1_1934_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1942_inst flow-through 
    process(BITSEL_u8_u1_1942_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1942_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1941_wire_constant = "& Convert_SLV_To_Hex_String(konst_1941_wire_constant) & " outputs:" & " BITSEL_u8_u1_1942_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1942_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1942_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1941_wire_constant, tmp_var);
      BITSEL_u8_u1_1942_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_194_inst flow-through 
    process(BITSEL_u8_u1_194_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_194_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_193_wire_constant = "& Convert_SLV_To_Hex_String(konst_193_wire_constant) & " outputs:" & " BITSEL_u8_u1_194_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_194_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_194_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_193_wire_constant, tmp_var);
      BITSEL_u8_u1_194_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1950_inst flow-through 
    process(BITSEL_u8_u1_1950_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1950_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1949_wire_constant = "& Convert_SLV_To_Hex_String(konst_1949_wire_constant) & " outputs:" & " BITSEL_u8_u1_1950_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1950_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1950_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1949_wire_constant, tmp_var);
      BITSEL_u8_u1_1950_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1958_inst flow-through 
    process(BITSEL_u8_u1_1958_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1958_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1957_wire_constant = "& Convert_SLV_To_Hex_String(konst_1957_wire_constant) & " outputs:" & " BITSEL_u8_u1_1958_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1958_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1958_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1957_wire_constant, tmp_var);
      BITSEL_u8_u1_1958_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1966_inst flow-through 
    process(BITSEL_u8_u1_1966_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1966_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1965_wire_constant = "& Convert_SLV_To_Hex_String(konst_1965_wire_constant) & " outputs:" & " BITSEL_u8_u1_1966_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1966_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1966_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1965_wire_constant, tmp_var);
      BITSEL_u8_u1_1966_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1974_inst flow-through 
    process(BITSEL_u8_u1_1974_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1974_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1973_wire_constant = "& Convert_SLV_To_Hex_String(konst_1973_wire_constant) & " outputs:" & " BITSEL_u8_u1_1974_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1974_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1974_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1973_wire_constant, tmp_var);
      BITSEL_u8_u1_1974_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1982_inst flow-through 
    process(BITSEL_u8_u1_1982_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1982_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1981_wire_constant = "& Convert_SLV_To_Hex_String(konst_1981_wire_constant) & " outputs:" & " BITSEL_u8_u1_1982_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1982_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1982_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1981_wire_constant, tmp_var);
      BITSEL_u8_u1_1982_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1990_inst flow-through 
    process(BITSEL_u8_u1_1990_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1990_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1989_wire_constant = "& Convert_SLV_To_Hex_String(konst_1989_wire_constant) & " outputs:" & " BITSEL_u8_u1_1990_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1990_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1990_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1989_wire_constant, tmp_var);
      BITSEL_u8_u1_1990_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_1998_inst flow-through 
    process(BITSEL_u8_u1_1998_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_1998_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_1997_wire_constant = "& Convert_SLV_To_Hex_String(konst_1997_wire_constant) & " outputs:" & " BITSEL_u8_u1_1998_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1998_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1998_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1997_wire_constant, tmp_var);
      BITSEL_u8_u1_1998_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_2006_inst flow-through 
    process(BITSEL_u8_u1_2006_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_2006_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_2005_wire_constant = "& Convert_SLV_To_Hex_String(konst_2005_wire_constant) & " outputs:" & " BITSEL_u8_u1_2006_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_2006_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_2006_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2005_wire_constant, tmp_var);
      BITSEL_u8_u1_2006_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_2014_inst flow-through 
    process(BITSEL_u8_u1_2014_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_2014_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_2013_wire_constant = "& Convert_SLV_To_Hex_String(konst_2013_wire_constant) & " outputs:" & " BITSEL_u8_u1_2014_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_2014_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_2014_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2013_wire_constant, tmp_var);
      BITSEL_u8_u1_2014_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_2022_inst flow-through 
    process(BITSEL_u8_u1_2022_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_2022_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_2021_wire_constant = "& Convert_SLV_To_Hex_String(konst_2021_wire_constant) & " outputs:" & " BITSEL_u8_u1_2022_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_2022_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_2022_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2021_wire_constant, tmp_var);
      BITSEL_u8_u1_2022_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_2030_inst flow-through 
    process(BITSEL_u8_u1_2030_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_2030_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_2029_wire_constant = "& Convert_SLV_To_Hex_String(konst_2029_wire_constant) & " outputs:" & " BITSEL_u8_u1_2030_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_2030_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_2030_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2029_wire_constant, tmp_var);
      BITSEL_u8_u1_2030_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_2038_inst flow-through 
    process(BITSEL_u8_u1_2038_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_2038_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_2037_wire_constant = "& Convert_SLV_To_Hex_String(konst_2037_wire_constant) & " outputs:" & " BITSEL_u8_u1_2038_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_2038_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_2038_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2037_wire_constant, tmp_var);
      BITSEL_u8_u1_2038_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_2046_inst flow-through 
    process(BITSEL_u8_u1_2046_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_2046_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_2045_wire_constant = "& Convert_SLV_To_Hex_String(konst_2045_wire_constant) & " outputs:" & " BITSEL_u8_u1_2046_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_2046_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_2046_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2045_wire_constant, tmp_var);
      BITSEL_u8_u1_2046_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_204_inst flow-through 
    process(BITSEL_u8_u1_204_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_204_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_203_wire_constant = "& Convert_SLV_To_Hex_String(konst_203_wire_constant) & " outputs:" & " BITSEL_u8_u1_204_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_204_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_204_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_203_wire_constant, tmp_var);
      BITSEL_u8_u1_204_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_2054_inst flow-through 
    process(BITSEL_u8_u1_2054_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_2054_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_2053_wire_constant = "& Convert_SLV_To_Hex_String(konst_2053_wire_constant) & " outputs:" & " BITSEL_u8_u1_2054_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_2054_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_2054_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2053_wire_constant, tmp_var);
      BITSEL_u8_u1_2054_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_2062_inst flow-through 
    process(BITSEL_u8_u1_2062_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_2062_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_2061_wire_constant = "& Convert_SLV_To_Hex_String(konst_2061_wire_constant) & " outputs:" & " BITSEL_u8_u1_2062_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_2062_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_2062_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2061_wire_constant, tmp_var);
      BITSEL_u8_u1_2062_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_2070_inst flow-through 
    process(BITSEL_u8_u1_2070_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_2070_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_2069_wire_constant = "& Convert_SLV_To_Hex_String(konst_2069_wire_constant) & " outputs:" & " BITSEL_u8_u1_2070_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_2070_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_2070_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2069_wire_constant, tmp_var);
      BITSEL_u8_u1_2070_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_2078_inst flow-through 
    process(BITSEL_u8_u1_2078_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_2078_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_2077_wire_constant = "& Convert_SLV_To_Hex_String(konst_2077_wire_constant) & " outputs:" & " BITSEL_u8_u1_2078_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_2078_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_2078_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2077_wire_constant, tmp_var);
      BITSEL_u8_u1_2078_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_2086_inst flow-through 
    process(BITSEL_u8_u1_2086_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_2086_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_2085_wire_constant = "& Convert_SLV_To_Hex_String(konst_2085_wire_constant) & " outputs:" & " BITSEL_u8_u1_2086_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_2086_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_2086_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2085_wire_constant, tmp_var);
      BITSEL_u8_u1_2086_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_2094_inst flow-through 
    process(BITSEL_u8_u1_2094_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_2094_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_2093_wire_constant = "& Convert_SLV_To_Hex_String(konst_2093_wire_constant) & " outputs:" & " BITSEL_u8_u1_2094_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_2094_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_2094_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2093_wire_constant, tmp_var);
      BITSEL_u8_u1_2094_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_2102_inst flow-through 
    process(BITSEL_u8_u1_2102_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_2102_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_2101_wire_constant = "& Convert_SLV_To_Hex_String(konst_2101_wire_constant) & " outputs:" & " BITSEL_u8_u1_2102_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_2102_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_2102_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2101_wire_constant, tmp_var);
      BITSEL_u8_u1_2102_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_2110_inst flow-through 
    process(BITSEL_u8_u1_2110_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_2110_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_2109_wire_constant = "& Convert_SLV_To_Hex_String(konst_2109_wire_constant) & " outputs:" & " BITSEL_u8_u1_2110_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_2110_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_2110_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2109_wire_constant, tmp_var);
      BITSEL_u8_u1_2110_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_2118_inst flow-through 
    process(BITSEL_u8_u1_2118_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_2118_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_2117_wire_constant = "& Convert_SLV_To_Hex_String(konst_2117_wire_constant) & " outputs:" & " BITSEL_u8_u1_2118_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_2118_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_2118_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2117_wire_constant, tmp_var);
      BITSEL_u8_u1_2118_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_2126_inst flow-through 
    process(BITSEL_u8_u1_2126_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_2126_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_2125_wire_constant = "& Convert_SLV_To_Hex_String(konst_2125_wire_constant) & " outputs:" & " BITSEL_u8_u1_2126_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_2126_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_2126_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2125_wire_constant, tmp_var);
      BITSEL_u8_u1_2126_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_2134_inst flow-through 
    process(BITSEL_u8_u1_2134_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_2134_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_2133_wire_constant = "& Convert_SLV_To_Hex_String(konst_2133_wire_constant) & " outputs:" & " BITSEL_u8_u1_2134_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_2134_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_2134_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2133_wire_constant, tmp_var);
      BITSEL_u8_u1_2134_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_2142_inst flow-through 
    process(BITSEL_u8_u1_2142_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_2142_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_2141_wire_constant = "& Convert_SLV_To_Hex_String(konst_2141_wire_constant) & " outputs:" & " BITSEL_u8_u1_2142_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_2142_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_2142_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2141_wire_constant, tmp_var);
      BITSEL_u8_u1_2142_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_214_inst flow-through 
    process(BITSEL_u8_u1_214_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_214_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_213_wire_constant = "& Convert_SLV_To_Hex_String(konst_213_wire_constant) & " outputs:" & " BITSEL_u8_u1_214_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_214_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_214_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_213_wire_constant, tmp_var);
      BITSEL_u8_u1_214_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_2150_inst flow-through 
    process(BITSEL_u8_u1_2150_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_2150_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_2149_wire_constant = "& Convert_SLV_To_Hex_String(konst_2149_wire_constant) & " outputs:" & " BITSEL_u8_u1_2150_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_2150_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_2150_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2149_wire_constant, tmp_var);
      BITSEL_u8_u1_2150_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_2158_inst flow-through 
    process(BITSEL_u8_u1_2158_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_2158_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_2157_wire_constant = "& Convert_SLV_To_Hex_String(konst_2157_wire_constant) & " outputs:" & " BITSEL_u8_u1_2158_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_2158_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_2158_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2157_wire_constant, tmp_var);
      BITSEL_u8_u1_2158_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_2166_inst flow-through 
    process(BITSEL_u8_u1_2166_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_2166_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_2165_wire_constant = "& Convert_SLV_To_Hex_String(konst_2165_wire_constant) & " outputs:" & " BITSEL_u8_u1_2166_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_2166_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_2166_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2165_wire_constant, tmp_var);
      BITSEL_u8_u1_2166_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_2174_inst flow-through 
    process(BITSEL_u8_u1_2174_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_2174_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_2173_wire_constant = "& Convert_SLV_To_Hex_String(konst_2173_wire_constant) & " outputs:" & " BITSEL_u8_u1_2174_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_2174_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_2174_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2173_wire_constant, tmp_var);
      BITSEL_u8_u1_2174_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_2182_inst flow-through 
    process(BITSEL_u8_u1_2182_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_2182_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_2181_wire_constant = "& Convert_SLV_To_Hex_String(konst_2181_wire_constant) & " outputs:" & " BITSEL_u8_u1_2182_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_2182_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_2182_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2181_wire_constant, tmp_var);
      BITSEL_u8_u1_2182_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_2190_inst flow-through 
    process(BITSEL_u8_u1_2190_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_2190_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_2189_wire_constant = "& Convert_SLV_To_Hex_String(konst_2189_wire_constant) & " outputs:" & " BITSEL_u8_u1_2190_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_2190_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_2190_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2189_wire_constant, tmp_var);
      BITSEL_u8_u1_2190_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_2198_inst flow-through 
    process(BITSEL_u8_u1_2198_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_2198_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_2197_wire_constant = "& Convert_SLV_To_Hex_String(konst_2197_wire_constant) & " outputs:" & " BITSEL_u8_u1_2198_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_2198_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_2198_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2197_wire_constant, tmp_var);
      BITSEL_u8_u1_2198_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_2206_inst flow-through 
    process(BITSEL_u8_u1_2206_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_2206_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_2205_wire_constant = "& Convert_SLV_To_Hex_String(konst_2205_wire_constant) & " outputs:" & " BITSEL_u8_u1_2206_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_2206_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_2206_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2205_wire_constant, tmp_var);
      BITSEL_u8_u1_2206_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_2214_inst flow-through 
    process(BITSEL_u8_u1_2214_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_2214_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_2213_wire_constant = "& Convert_SLV_To_Hex_String(konst_2213_wire_constant) & " outputs:" & " BITSEL_u8_u1_2214_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_2214_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_2214_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2213_wire_constant, tmp_var);
      BITSEL_u8_u1_2214_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_2222_inst flow-through 
    process(BITSEL_u8_u1_2222_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_2222_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_2221_wire_constant = "& Convert_SLV_To_Hex_String(konst_2221_wire_constant) & " outputs:" & " BITSEL_u8_u1_2222_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_2222_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_2222_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2221_wire_constant, tmp_var);
      BITSEL_u8_u1_2222_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_2230_inst flow-through 
    process(BITSEL_u8_u1_2230_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_2230_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_2229_wire_constant = "& Convert_SLV_To_Hex_String(konst_2229_wire_constant) & " outputs:" & " BITSEL_u8_u1_2230_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_2230_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_2230_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2229_wire_constant, tmp_var);
      BITSEL_u8_u1_2230_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_2238_inst flow-through 
    process(BITSEL_u8_u1_2238_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_2238_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_2237_wire_constant = "& Convert_SLV_To_Hex_String(konst_2237_wire_constant) & " outputs:" & " BITSEL_u8_u1_2238_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_2238_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_2238_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2237_wire_constant, tmp_var);
      BITSEL_u8_u1_2238_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_2246_inst flow-through 
    process(BITSEL_u8_u1_2246_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_2246_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_2245_wire_constant = "& Convert_SLV_To_Hex_String(konst_2245_wire_constant) & " outputs:" & " BITSEL_u8_u1_2246_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_2246_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_2246_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2245_wire_constant, tmp_var);
      BITSEL_u8_u1_2246_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_224_inst flow-through 
    process(BITSEL_u8_u1_224_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_224_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_223_wire_constant = "& Convert_SLV_To_Hex_String(konst_223_wire_constant) & " outputs:" & " BITSEL_u8_u1_224_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_224_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_224_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_223_wire_constant, tmp_var);
      BITSEL_u8_u1_224_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_2254_inst flow-through 
    process(BITSEL_u8_u1_2254_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_2254_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_2253_wire_constant = "& Convert_SLV_To_Hex_String(konst_2253_wire_constant) & " outputs:" & " BITSEL_u8_u1_2254_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_2254_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_2254_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2253_wire_constant, tmp_var);
      BITSEL_u8_u1_2254_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_2262_inst flow-through 
    process(BITSEL_u8_u1_2262_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_2262_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_2261_wire_constant = "& Convert_SLV_To_Hex_String(konst_2261_wire_constant) & " outputs:" & " BITSEL_u8_u1_2262_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_2262_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_2262_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2261_wire_constant, tmp_var);
      BITSEL_u8_u1_2262_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_2270_inst flow-through 
    process(BITSEL_u8_u1_2270_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_2270_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_2269_wire_constant = "& Convert_SLV_To_Hex_String(konst_2269_wire_constant) & " outputs:" & " BITSEL_u8_u1_2270_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_2270_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_2270_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2269_wire_constant, tmp_var);
      BITSEL_u8_u1_2270_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_2278_inst flow-through 
    process(BITSEL_u8_u1_2278_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_2278_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_2277_wire_constant = "& Convert_SLV_To_Hex_String(konst_2277_wire_constant) & " outputs:" & " BITSEL_u8_u1_2278_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_2278_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_2278_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2277_wire_constant, tmp_var);
      BITSEL_u8_u1_2278_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_2286_inst flow-through 
    process(BITSEL_u8_u1_2286_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_2286_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_2285_wire_constant = "& Convert_SLV_To_Hex_String(konst_2285_wire_constant) & " outputs:" & " BITSEL_u8_u1_2286_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_2286_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_2286_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2285_wire_constant, tmp_var);
      BITSEL_u8_u1_2286_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_2294_inst flow-through 
    process(BITSEL_u8_u1_2294_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_2294_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_2293_wire_constant = "& Convert_SLV_To_Hex_String(konst_2293_wire_constant) & " outputs:" & " BITSEL_u8_u1_2294_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_2294_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_2294_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2293_wire_constant, tmp_var);
      BITSEL_u8_u1_2294_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_2302_inst flow-through 
    process(BITSEL_u8_u1_2302_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_2302_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_2301_wire_constant = "& Convert_SLV_To_Hex_String(konst_2301_wire_constant) & " outputs:" & " BITSEL_u8_u1_2302_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_2302_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_2302_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2301_wire_constant, tmp_var);
      BITSEL_u8_u1_2302_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_234_inst flow-through 
    process(BITSEL_u8_u1_234_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_234_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_233_wire_constant = "& Convert_SLV_To_Hex_String(konst_233_wire_constant) & " outputs:" & " BITSEL_u8_u1_234_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_234_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_234_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_233_wire_constant, tmp_var);
      BITSEL_u8_u1_234_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_244_inst flow-through 
    process(BITSEL_u8_u1_244_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_244_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_243_wire_constant = "& Convert_SLV_To_Hex_String(konst_243_wire_constant) & " outputs:" & " BITSEL_u8_u1_244_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_244_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_244_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_243_wire_constant, tmp_var);
      BITSEL_u8_u1_244_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_24_inst flow-through 
    process(BITSEL_u8_u1_24_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_24_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_23_wire_constant = "& Convert_SLV_To_Hex_String(konst_23_wire_constant) & " outputs:" & " BITSEL_u8_u1_24_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_24_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_24_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_23_wire_constant, tmp_var);
      BITSEL_u8_u1_24_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_254_inst flow-through 
    process(BITSEL_u8_u1_254_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_254_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_253_wire_constant = "& Convert_SLV_To_Hex_String(konst_253_wire_constant) & " outputs:" & " BITSEL_u8_u1_254_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_254_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_254_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_253_wire_constant, tmp_var);
      BITSEL_u8_u1_254_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_264_inst flow-through 
    process(BITSEL_u8_u1_264_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_264_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_263_wire_constant = "& Convert_SLV_To_Hex_String(konst_263_wire_constant) & " outputs:" & " BITSEL_u8_u1_264_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_264_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_264_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_263_wire_constant, tmp_var);
      BITSEL_u8_u1_264_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_274_inst flow-through 
    process(BITSEL_u8_u1_274_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_274_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_273_wire_constant = "& Convert_SLV_To_Hex_String(konst_273_wire_constant) & " outputs:" & " BITSEL_u8_u1_274_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_274_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_274_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_273_wire_constant, tmp_var);
      BITSEL_u8_u1_274_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_284_inst flow-through 
    process(BITSEL_u8_u1_284_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_284_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_283_wire_constant = "& Convert_SLV_To_Hex_String(konst_283_wire_constant) & " outputs:" & " BITSEL_u8_u1_284_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_284_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_284_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_283_wire_constant, tmp_var);
      BITSEL_u8_u1_284_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_294_inst flow-through 
    process(BITSEL_u8_u1_294_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_294_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_293_wire_constant = "& Convert_SLV_To_Hex_String(konst_293_wire_constant) & " outputs:" & " BITSEL_u8_u1_294_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_294_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_294_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_293_wire_constant, tmp_var);
      BITSEL_u8_u1_294_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_304_inst flow-through 
    process(BITSEL_u8_u1_304_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_304_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_303_wire_constant = "& Convert_SLV_To_Hex_String(konst_303_wire_constant) & " outputs:" & " BITSEL_u8_u1_304_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_304_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_304_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_303_wire_constant, tmp_var);
      BITSEL_u8_u1_304_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_314_inst flow-through 
    process(BITSEL_u8_u1_314_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_314_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_313_wire_constant = "& Convert_SLV_To_Hex_String(konst_313_wire_constant) & " outputs:" & " BITSEL_u8_u1_314_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_314_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_314_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_313_wire_constant, tmp_var);
      BITSEL_u8_u1_314_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_324_inst flow-through 
    process(BITSEL_u8_u1_324_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_324_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_323_wire_constant = "& Convert_SLV_To_Hex_String(konst_323_wire_constant) & " outputs:" & " BITSEL_u8_u1_324_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_324_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_324_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_323_wire_constant, tmp_var);
      BITSEL_u8_u1_324_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_334_inst flow-through 
    process(BITSEL_u8_u1_334_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_334_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_333_wire_constant = "& Convert_SLV_To_Hex_String(konst_333_wire_constant) & " outputs:" & " BITSEL_u8_u1_334_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_334_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_334_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_333_wire_constant, tmp_var);
      BITSEL_u8_u1_334_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_344_inst flow-through 
    process(BITSEL_u8_u1_344_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_344_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_343_wire_constant = "& Convert_SLV_To_Hex_String(konst_343_wire_constant) & " outputs:" & " BITSEL_u8_u1_344_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_344_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_344_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_343_wire_constant, tmp_var);
      BITSEL_u8_u1_344_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_34_inst flow-through 
    process(BITSEL_u8_u1_34_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_34_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_33_wire_constant = "& Convert_SLV_To_Hex_String(konst_33_wire_constant) & " outputs:" & " BITSEL_u8_u1_34_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_34_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_34_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_33_wire_constant, tmp_var);
      BITSEL_u8_u1_34_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_354_inst flow-through 
    process(BITSEL_u8_u1_354_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_354_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_353_wire_constant = "& Convert_SLV_To_Hex_String(konst_353_wire_constant) & " outputs:" & " BITSEL_u8_u1_354_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_354_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_354_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_353_wire_constant, tmp_var);
      BITSEL_u8_u1_354_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_364_inst flow-through 
    process(BITSEL_u8_u1_364_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_364_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_363_wire_constant = "& Convert_SLV_To_Hex_String(konst_363_wire_constant) & " outputs:" & " BITSEL_u8_u1_364_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_364_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_364_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_363_wire_constant, tmp_var);
      BITSEL_u8_u1_364_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_374_inst flow-through 
    process(BITSEL_u8_u1_374_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_374_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_373_wire_constant = "& Convert_SLV_To_Hex_String(konst_373_wire_constant) & " outputs:" & " BITSEL_u8_u1_374_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_374_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_374_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_373_wire_constant, tmp_var);
      BITSEL_u8_u1_374_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_384_inst flow-through 
    process(BITSEL_u8_u1_384_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_384_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_383_wire_constant = "& Convert_SLV_To_Hex_String(konst_383_wire_constant) & " outputs:" & " BITSEL_u8_u1_384_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_384_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_384_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_383_wire_constant, tmp_var);
      BITSEL_u8_u1_384_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_394_inst flow-through 
    process(BITSEL_u8_u1_394_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_394_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_393_wire_constant = "& Convert_SLV_To_Hex_String(konst_393_wire_constant) & " outputs:" & " BITSEL_u8_u1_394_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_394_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_394_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_393_wire_constant, tmp_var);
      BITSEL_u8_u1_394_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_404_inst flow-through 
    process(BITSEL_u8_u1_404_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_404_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_403_wire_constant = "& Convert_SLV_To_Hex_String(konst_403_wire_constant) & " outputs:" & " BITSEL_u8_u1_404_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_404_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_404_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_403_wire_constant, tmp_var);
      BITSEL_u8_u1_404_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_414_inst flow-through 
    process(BITSEL_u8_u1_414_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_414_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_413_wire_constant = "& Convert_SLV_To_Hex_String(konst_413_wire_constant) & " outputs:" & " BITSEL_u8_u1_414_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_414_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_414_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_413_wire_constant, tmp_var);
      BITSEL_u8_u1_414_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_424_inst flow-through 
    process(BITSEL_u8_u1_424_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_424_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_423_wire_constant = "& Convert_SLV_To_Hex_String(konst_423_wire_constant) & " outputs:" & " BITSEL_u8_u1_424_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_424_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_424_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_423_wire_constant, tmp_var);
      BITSEL_u8_u1_424_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_434_inst flow-through 
    process(BITSEL_u8_u1_434_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_434_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_433_wire_constant = "& Convert_SLV_To_Hex_String(konst_433_wire_constant) & " outputs:" & " BITSEL_u8_u1_434_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_434_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_434_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_433_wire_constant, tmp_var);
      BITSEL_u8_u1_434_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_444_inst flow-through 
    process(BITSEL_u8_u1_444_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_444_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_443_wire_constant = "& Convert_SLV_To_Hex_String(konst_443_wire_constant) & " outputs:" & " BITSEL_u8_u1_444_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_444_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_444_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_443_wire_constant, tmp_var);
      BITSEL_u8_u1_444_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_44_inst flow-through 
    process(BITSEL_u8_u1_44_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_44_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_43_wire_constant = "& Convert_SLV_To_Hex_String(konst_43_wire_constant) & " outputs:" & " BITSEL_u8_u1_44_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_44_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_44_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_43_wire_constant, tmp_var);
      BITSEL_u8_u1_44_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_454_inst flow-through 
    process(BITSEL_u8_u1_454_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_454_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_453_wire_constant = "& Convert_SLV_To_Hex_String(konst_453_wire_constant) & " outputs:" & " BITSEL_u8_u1_454_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_454_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_454_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_453_wire_constant, tmp_var);
      BITSEL_u8_u1_454_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_464_inst flow-through 
    process(BITSEL_u8_u1_464_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_464_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_463_wire_constant = "& Convert_SLV_To_Hex_String(konst_463_wire_constant) & " outputs:" & " BITSEL_u8_u1_464_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_464_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_464_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_463_wire_constant, tmp_var);
      BITSEL_u8_u1_464_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_474_inst flow-through 
    process(BITSEL_u8_u1_474_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_474_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_473_wire_constant = "& Convert_SLV_To_Hex_String(konst_473_wire_constant) & " outputs:" & " BITSEL_u8_u1_474_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_474_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_474_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_473_wire_constant, tmp_var);
      BITSEL_u8_u1_474_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_484_inst flow-through 
    process(BITSEL_u8_u1_484_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_484_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_483_wire_constant = "& Convert_SLV_To_Hex_String(konst_483_wire_constant) & " outputs:" & " BITSEL_u8_u1_484_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_484_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_484_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_483_wire_constant, tmp_var);
      BITSEL_u8_u1_484_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_494_inst flow-through 
    process(BITSEL_u8_u1_494_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_494_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_493_wire_constant = "& Convert_SLV_To_Hex_String(konst_493_wire_constant) & " outputs:" & " BITSEL_u8_u1_494_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_494_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_494_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_493_wire_constant, tmp_var);
      BITSEL_u8_u1_494_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_504_inst flow-through 
    process(BITSEL_u8_u1_504_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_504_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_503_wire_constant = "& Convert_SLV_To_Hex_String(konst_503_wire_constant) & " outputs:" & " BITSEL_u8_u1_504_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_504_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_504_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_503_wire_constant, tmp_var);
      BITSEL_u8_u1_504_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_514_inst flow-through 
    process(BITSEL_u8_u1_514_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_514_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_513_wire_constant = "& Convert_SLV_To_Hex_String(konst_513_wire_constant) & " outputs:" & " BITSEL_u8_u1_514_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_514_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_514_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_513_wire_constant, tmp_var);
      BITSEL_u8_u1_514_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_524_inst flow-through 
    process(BITSEL_u8_u1_524_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_524_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_523_wire_constant = "& Convert_SLV_To_Hex_String(konst_523_wire_constant) & " outputs:" & " BITSEL_u8_u1_524_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_524_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_524_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_523_wire_constant, tmp_var);
      BITSEL_u8_u1_524_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_534_inst flow-through 
    process(BITSEL_u8_u1_534_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_534_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_533_wire_constant = "& Convert_SLV_To_Hex_String(konst_533_wire_constant) & " outputs:" & " BITSEL_u8_u1_534_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_534_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_534_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_533_wire_constant, tmp_var);
      BITSEL_u8_u1_534_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_544_inst flow-through 
    process(BITSEL_u8_u1_544_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_544_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_543_wire_constant = "& Convert_SLV_To_Hex_String(konst_543_wire_constant) & " outputs:" & " BITSEL_u8_u1_544_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_544_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_544_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_543_wire_constant, tmp_var);
      BITSEL_u8_u1_544_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_54_inst flow-through 
    process(BITSEL_u8_u1_54_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_54_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_53_wire_constant = "& Convert_SLV_To_Hex_String(konst_53_wire_constant) & " outputs:" & " BITSEL_u8_u1_54_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_54_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_54_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_53_wire_constant, tmp_var);
      BITSEL_u8_u1_54_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_554_inst flow-through 
    process(BITSEL_u8_u1_554_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_554_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_553_wire_constant = "& Convert_SLV_To_Hex_String(konst_553_wire_constant) & " outputs:" & " BITSEL_u8_u1_554_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_554_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_554_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_553_wire_constant, tmp_var);
      BITSEL_u8_u1_554_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_564_inst flow-through 
    process(BITSEL_u8_u1_564_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_564_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_563_wire_constant = "& Convert_SLV_To_Hex_String(konst_563_wire_constant) & " outputs:" & " BITSEL_u8_u1_564_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_564_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_564_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_563_wire_constant, tmp_var);
      BITSEL_u8_u1_564_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_574_inst flow-through 
    process(BITSEL_u8_u1_574_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_574_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_573_wire_constant = "& Convert_SLV_To_Hex_String(konst_573_wire_constant) & " outputs:" & " BITSEL_u8_u1_574_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_574_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_574_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_573_wire_constant, tmp_var);
      BITSEL_u8_u1_574_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_584_inst flow-through 
    process(BITSEL_u8_u1_584_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_584_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_583_wire_constant = "& Convert_SLV_To_Hex_String(konst_583_wire_constant) & " outputs:" & " BITSEL_u8_u1_584_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_584_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_584_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_583_wire_constant, tmp_var);
      BITSEL_u8_u1_584_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_594_inst flow-through 
    process(BITSEL_u8_u1_594_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_594_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_593_wire_constant = "& Convert_SLV_To_Hex_String(konst_593_wire_constant) & " outputs:" & " BITSEL_u8_u1_594_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_594_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_594_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_593_wire_constant, tmp_var);
      BITSEL_u8_u1_594_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_604_inst flow-through 
    process(BITSEL_u8_u1_604_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_604_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_603_wire_constant = "& Convert_SLV_To_Hex_String(konst_603_wire_constant) & " outputs:" & " BITSEL_u8_u1_604_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_604_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_604_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_603_wire_constant, tmp_var);
      BITSEL_u8_u1_604_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_614_inst flow-through 
    process(BITSEL_u8_u1_614_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_614_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_613_wire_constant = "& Convert_SLV_To_Hex_String(konst_613_wire_constant) & " outputs:" & " BITSEL_u8_u1_614_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_614_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_614_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_613_wire_constant, tmp_var);
      BITSEL_u8_u1_614_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_624_inst flow-through 
    process(BITSEL_u8_u1_624_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_624_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_623_wire_constant = "& Convert_SLV_To_Hex_String(konst_623_wire_constant) & " outputs:" & " BITSEL_u8_u1_624_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_624_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_624_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_623_wire_constant, tmp_var);
      BITSEL_u8_u1_624_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_634_inst flow-through 
    process(BITSEL_u8_u1_634_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_634_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_633_wire_constant = "& Convert_SLV_To_Hex_String(konst_633_wire_constant) & " outputs:" & " BITSEL_u8_u1_634_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_634_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_634_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_633_wire_constant, tmp_var);
      BITSEL_u8_u1_634_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_644_inst flow-through 
    process(BITSEL_u8_u1_644_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_644_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_643_wire_constant = "& Convert_SLV_To_Hex_String(konst_643_wire_constant) & " outputs:" & " BITSEL_u8_u1_644_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_644_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_644_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_643_wire_constant, tmp_var);
      BITSEL_u8_u1_644_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_64_inst flow-through 
    process(BITSEL_u8_u1_64_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_64_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_63_wire_constant = "& Convert_SLV_To_Hex_String(konst_63_wire_constant) & " outputs:" & " BITSEL_u8_u1_64_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_64_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_64_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_63_wire_constant, tmp_var);
      BITSEL_u8_u1_64_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_654_inst flow-through 
    process(BITSEL_u8_u1_654_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_654_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_653_wire_constant = "& Convert_SLV_To_Hex_String(konst_653_wire_constant) & " outputs:" & " BITSEL_u8_u1_654_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_654_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_654_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_653_wire_constant, tmp_var);
      BITSEL_u8_u1_654_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_664_inst flow-through 
    process(BITSEL_u8_u1_664_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_664_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_663_wire_constant = "& Convert_SLV_To_Hex_String(konst_663_wire_constant) & " outputs:" & " BITSEL_u8_u1_664_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_664_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_664_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_663_wire_constant, tmp_var);
      BITSEL_u8_u1_664_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_674_inst flow-through 
    process(BITSEL_u8_u1_674_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_674_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_673_wire_constant = "& Convert_SLV_To_Hex_String(konst_673_wire_constant) & " outputs:" & " BITSEL_u8_u1_674_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_674_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_674_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_673_wire_constant, tmp_var);
      BITSEL_u8_u1_674_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_684_inst flow-through 
    process(BITSEL_u8_u1_684_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_684_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_683_wire_constant = "& Convert_SLV_To_Hex_String(konst_683_wire_constant) & " outputs:" & " BITSEL_u8_u1_684_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_684_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_684_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_683_wire_constant, tmp_var);
      BITSEL_u8_u1_684_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_694_inst flow-through 
    process(BITSEL_u8_u1_694_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_694_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_693_wire_constant = "& Convert_SLV_To_Hex_String(konst_693_wire_constant) & " outputs:" & " BITSEL_u8_u1_694_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_694_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_694_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_693_wire_constant, tmp_var);
      BITSEL_u8_u1_694_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_704_inst flow-through 
    process(BITSEL_u8_u1_704_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_704_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_703_wire_constant = "& Convert_SLV_To_Hex_String(konst_703_wire_constant) & " outputs:" & " BITSEL_u8_u1_704_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_704_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_704_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_703_wire_constant, tmp_var);
      BITSEL_u8_u1_704_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_714_inst flow-through 
    process(BITSEL_u8_u1_714_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_714_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_713_wire_constant = "& Convert_SLV_To_Hex_String(konst_713_wire_constant) & " outputs:" & " BITSEL_u8_u1_714_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_714_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_714_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_713_wire_constant, tmp_var);
      BITSEL_u8_u1_714_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_724_inst flow-through 
    process(BITSEL_u8_u1_724_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_724_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_723_wire_constant = "& Convert_SLV_To_Hex_String(konst_723_wire_constant) & " outputs:" & " BITSEL_u8_u1_724_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_724_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_724_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_723_wire_constant, tmp_var);
      BITSEL_u8_u1_724_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_734_inst flow-through 
    process(BITSEL_u8_u1_734_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_734_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_733_wire_constant = "& Convert_SLV_To_Hex_String(konst_733_wire_constant) & " outputs:" & " BITSEL_u8_u1_734_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_734_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_734_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_733_wire_constant, tmp_var);
      BITSEL_u8_u1_734_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_744_inst flow-through 
    process(BITSEL_u8_u1_744_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_744_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_743_wire_constant = "& Convert_SLV_To_Hex_String(konst_743_wire_constant) & " outputs:" & " BITSEL_u8_u1_744_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_744_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_744_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_743_wire_constant, tmp_var);
      BITSEL_u8_u1_744_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_74_inst flow-through 
    process(BITSEL_u8_u1_74_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_74_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_73_wire_constant = "& Convert_SLV_To_Hex_String(konst_73_wire_constant) & " outputs:" & " BITSEL_u8_u1_74_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_74_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_74_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_73_wire_constant, tmp_var);
      BITSEL_u8_u1_74_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_754_inst flow-through 
    process(BITSEL_u8_u1_754_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_754_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_753_wire_constant = "& Convert_SLV_To_Hex_String(konst_753_wire_constant) & " outputs:" & " BITSEL_u8_u1_754_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_754_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_754_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_753_wire_constant, tmp_var);
      BITSEL_u8_u1_754_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_764_inst flow-through 
    process(BITSEL_u8_u1_764_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_764_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_763_wire_constant = "& Convert_SLV_To_Hex_String(konst_763_wire_constant) & " outputs:" & " BITSEL_u8_u1_764_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_764_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_764_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_763_wire_constant, tmp_var);
      BITSEL_u8_u1_764_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_774_inst flow-through 
    process(BITSEL_u8_u1_774_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_774_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_773_wire_constant = "& Convert_SLV_To_Hex_String(konst_773_wire_constant) & " outputs:" & " BITSEL_u8_u1_774_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_774_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_774_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_773_wire_constant, tmp_var);
      BITSEL_u8_u1_774_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_784_inst flow-through 
    process(BITSEL_u8_u1_784_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_784_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_783_wire_constant = "& Convert_SLV_To_Hex_String(konst_783_wire_constant) & " outputs:" & " BITSEL_u8_u1_784_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_784_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_784_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_783_wire_constant, tmp_var);
      BITSEL_u8_u1_784_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_794_inst flow-through 
    process(BITSEL_u8_u1_794_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_794_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_793_wire_constant = "& Convert_SLV_To_Hex_String(konst_793_wire_constant) & " outputs:" & " BITSEL_u8_u1_794_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_794_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_794_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_793_wire_constant, tmp_var);
      BITSEL_u8_u1_794_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_804_inst flow-through 
    process(BITSEL_u8_u1_804_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_804_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_803_wire_constant = "& Convert_SLV_To_Hex_String(konst_803_wire_constant) & " outputs:" & " BITSEL_u8_u1_804_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_804_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_804_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_803_wire_constant, tmp_var);
      BITSEL_u8_u1_804_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_814_inst flow-through 
    process(BITSEL_u8_u1_814_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_814_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_813_wire_constant = "& Convert_SLV_To_Hex_String(konst_813_wire_constant) & " outputs:" & " BITSEL_u8_u1_814_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_814_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_814_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_813_wire_constant, tmp_var);
      BITSEL_u8_u1_814_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_824_inst flow-through 
    process(BITSEL_u8_u1_824_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_824_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_823_wire_constant = "& Convert_SLV_To_Hex_String(konst_823_wire_constant) & " outputs:" & " BITSEL_u8_u1_824_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_824_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_824_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_823_wire_constant, tmp_var);
      BITSEL_u8_u1_824_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_834_inst flow-through 
    process(BITSEL_u8_u1_834_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_834_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_833_wire_constant = "& Convert_SLV_To_Hex_String(konst_833_wire_constant) & " outputs:" & " BITSEL_u8_u1_834_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_834_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_834_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_833_wire_constant, tmp_var);
      BITSEL_u8_u1_834_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_844_inst flow-through 
    process(BITSEL_u8_u1_844_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_844_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_843_wire_constant = "& Convert_SLV_To_Hex_String(konst_843_wire_constant) & " outputs:" & " BITSEL_u8_u1_844_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_844_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_844_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_843_wire_constant, tmp_var);
      BITSEL_u8_u1_844_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_84_inst flow-through 
    process(BITSEL_u8_u1_84_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_84_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_83_wire_constant = "& Convert_SLV_To_Hex_String(konst_83_wire_constant) & " outputs:" & " BITSEL_u8_u1_84_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_84_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_84_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_83_wire_constant, tmp_var);
      BITSEL_u8_u1_84_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_854_inst flow-through 
    process(BITSEL_u8_u1_854_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_854_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_853_wire_constant = "& Convert_SLV_To_Hex_String(konst_853_wire_constant) & " outputs:" & " BITSEL_u8_u1_854_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_854_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_854_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_853_wire_constant, tmp_var);
      BITSEL_u8_u1_854_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_864_inst flow-through 
    process(BITSEL_u8_u1_864_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_864_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_863_wire_constant = "& Convert_SLV_To_Hex_String(konst_863_wire_constant) & " outputs:" & " BITSEL_u8_u1_864_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_864_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_864_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_863_wire_constant, tmp_var);
      BITSEL_u8_u1_864_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_874_inst flow-through 
    process(BITSEL_u8_u1_874_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_874_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_873_wire_constant = "& Convert_SLV_To_Hex_String(konst_873_wire_constant) & " outputs:" & " BITSEL_u8_u1_874_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_874_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_874_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_873_wire_constant, tmp_var);
      BITSEL_u8_u1_874_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_884_inst flow-through 
    process(BITSEL_u8_u1_884_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_884_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_883_wire_constant = "& Convert_SLV_To_Hex_String(konst_883_wire_constant) & " outputs:" & " BITSEL_u8_u1_884_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_884_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_884_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_883_wire_constant, tmp_var);
      BITSEL_u8_u1_884_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_894_inst flow-through 
    process(BITSEL_u8_u1_894_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_894_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_893_wire_constant = "& Convert_SLV_To_Hex_String(konst_893_wire_constant) & " outputs:" & " BITSEL_u8_u1_894_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_894_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_894_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_893_wire_constant, tmp_var);
      BITSEL_u8_u1_894_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_904_inst flow-through 
    process(BITSEL_u8_u1_904_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_904_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_903_wire_constant = "& Convert_SLV_To_Hex_String(konst_903_wire_constant) & " outputs:" & " BITSEL_u8_u1_904_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_904_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_904_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_903_wire_constant, tmp_var);
      BITSEL_u8_u1_904_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_914_inst flow-through 
    process(BITSEL_u8_u1_914_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_914_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_913_wire_constant = "& Convert_SLV_To_Hex_String(konst_913_wire_constant) & " outputs:" & " BITSEL_u8_u1_914_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_914_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_914_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_913_wire_constant, tmp_var);
      BITSEL_u8_u1_914_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_924_inst flow-through 
    process(BITSEL_u8_u1_924_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_924_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_923_wire_constant = "& Convert_SLV_To_Hex_String(konst_923_wire_constant) & " outputs:" & " BITSEL_u8_u1_924_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_924_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_924_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_923_wire_constant, tmp_var);
      BITSEL_u8_u1_924_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_934_inst flow-through 
    process(BITSEL_u8_u1_934_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_934_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_933_wire_constant = "& Convert_SLV_To_Hex_String(konst_933_wire_constant) & " outputs:" & " BITSEL_u8_u1_934_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_934_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_934_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_933_wire_constant, tmp_var);
      BITSEL_u8_u1_934_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_944_inst flow-through 
    process(BITSEL_u8_u1_944_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_944_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_943_wire_constant = "& Convert_SLV_To_Hex_String(konst_943_wire_constant) & " outputs:" & " BITSEL_u8_u1_944_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_944_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_944_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_943_wire_constant, tmp_var);
      BITSEL_u8_u1_944_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_94_inst flow-through 
    process(BITSEL_u8_u1_94_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_94_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_93_wire_constant = "& Convert_SLV_To_Hex_String(konst_93_wire_constant) & " outputs:" & " BITSEL_u8_u1_94_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_94_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_94_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_93_wire_constant, tmp_var);
      BITSEL_u8_u1_94_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_954_inst flow-through 
    process(BITSEL_u8_u1_954_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_954_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_953_wire_constant = "& Convert_SLV_To_Hex_String(konst_953_wire_constant) & " outputs:" & " BITSEL_u8_u1_954_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_954_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_954_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_953_wire_constant, tmp_var);
      BITSEL_u8_u1_954_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_964_inst flow-through 
    process(BITSEL_u8_u1_964_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_964_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_963_wire_constant = "& Convert_SLV_To_Hex_String(konst_963_wire_constant) & " outputs:" & " BITSEL_u8_u1_964_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_964_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_964_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_963_wire_constant, tmp_var);
      BITSEL_u8_u1_964_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_974_inst flow-through 
    process(BITSEL_u8_u1_974_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_974_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_973_wire_constant = "& Convert_SLV_To_Hex_String(konst_973_wire_constant) & " outputs:" & " BITSEL_u8_u1_974_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_974_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_974_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_973_wire_constant, tmp_var);
      BITSEL_u8_u1_974_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_984_inst flow-through 
    process(BITSEL_u8_u1_984_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_984_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_983_wire_constant = "& Convert_SLV_To_Hex_String(konst_983_wire_constant) & " outputs:" & " BITSEL_u8_u1_984_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_984_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_984_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_983_wire_constant, tmp_var);
      BITSEL_u8_u1_984_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_994_inst flow-through 
    process(BITSEL_u8_u1_994_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_1:DP:BITSEL_u8_u1_994_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_993_wire_constant = "& Convert_SLV_To_Hex_String(konst_993_wire_constant) & " outputs:" & " BITSEL_u8_u1_994_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_994_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_994_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_993_wire_constant, tmp_var);
      BITSEL_u8_u1_994_wire <= tmp_var; -- 
    end process;
    -- 
  end Block; -- data_path
  -- 
end Inv_Sbox_1_Volatile_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library GhdlLink;
use GhdlLink.LogUtilities.all;
library work;
use work.ahir_system_global_package.all;
entity Inv_Sbox_2_Volatile is -- 
  port ( -- 
    clk, reset: in std_logic; 
    s_in : in  std_logic_vector(7 downto 0);
    s_out : out  std_logic_vector(7 downto 0)-- 
  );
  -- 
end entity Inv_Sbox_2_Volatile;
architecture Inv_Sbox_2_Volatile_arch of Inv_Sbox_2_Volatile is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector(8-1 downto 0);
  signal default_zero_sig: std_logic;
  -- input port buffer signals
  signal s_in_buffer :  std_logic_vector(7 downto 0);
  -- output port buffer signals
  signal s_out_buffer :  std_logic_vector(7 downto 0);
  -- volatile/operator module components. 
  signal global_clock_cycle_count: integer := 0;
  -- 
begin --  
  ---------------------------------------------------------- 
  process(clk)  
  begin -- 
    if(clk'event and clk = '1') then -- 
      if(reset = '1') then -- 
        global_clock_cycle_count <= 0; --
      else -- 
        global_clock_cycle_count <= global_clock_cycle_count + 1; -- 
      end if; --
    end if; --
  end process;
  ---------------------------------------------------------- 
  -- input handling ------------------------------------------------
  s_in_buffer <= s_in;
  -- output handling  -------------------------------------------------------
  s_out <= s_out_buffer;
  -- the control path --------------------------------------------------
  default_zero_sig <= '0';
  -- volatile module, no control path
  -- the data path
  data_path: Block -- 
    signal BITSEL_u8_u1_2314_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2324_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2334_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2344_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2354_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2364_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2374_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2384_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2394_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2404_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2414_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2424_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2434_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2444_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2454_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2464_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2474_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2484_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2494_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2504_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2514_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2524_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2534_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2544_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2554_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2564_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2574_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2584_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2594_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2604_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2614_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2624_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2634_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2644_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2654_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2664_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2674_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2684_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2694_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2704_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2714_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2724_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2734_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2744_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2754_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2764_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2774_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2784_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2794_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2804_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2814_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2824_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2834_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2844_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2854_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2864_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2874_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2884_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2894_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2904_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2914_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2924_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2934_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2944_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2954_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2964_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2974_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2984_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2994_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3004_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3014_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3024_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3034_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3044_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3054_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3064_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3074_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3084_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3094_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3104_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3114_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3124_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3134_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3144_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3154_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3164_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3174_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3184_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3194_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3204_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3214_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3224_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3234_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3244_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3254_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3264_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3274_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3284_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3294_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3304_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3314_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3324_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3334_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3344_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3354_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3364_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3374_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3384_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3394_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3404_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3414_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3424_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3434_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3444_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3454_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3464_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3474_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3484_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3494_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3504_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3514_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3524_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3534_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3544_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3554_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3564_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3574_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3584_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3594_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3602_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3610_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3618_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3626_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3634_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3642_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3650_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3658_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3666_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3674_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3682_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3690_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3698_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3706_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3714_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3722_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3730_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3738_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3746_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3754_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3762_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3770_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3778_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3786_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3794_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3802_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3810_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3818_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3826_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3834_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3842_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3850_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3858_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3866_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3874_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3882_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3890_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3898_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3906_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3914_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3922_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3930_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3938_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3946_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3954_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3962_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3970_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3978_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3986_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3994_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4002_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4010_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4018_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4026_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4034_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4042_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4050_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4058_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4066_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4074_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4082_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4090_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4098_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4106_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4114_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4122_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4130_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4138_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4146_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4154_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4162_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4170_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4178_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4186_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4194_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4202_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4210_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4218_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4226_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4234_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4242_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4250_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4258_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4266_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4274_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4282_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4290_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4298_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4306_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4314_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4322_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4330_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4338_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4346_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4354_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4362_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4370_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4378_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4386_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4394_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4402_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4410_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4418_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4426_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4434_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4442_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4450_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4458_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4466_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4474_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4482_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4490_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4498_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4506_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4514_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4522_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4530_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4538_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4546_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4554_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4562_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4570_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4578_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4586_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4594_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4602_wire : std_logic_vector(0 downto 0);
    signal IMA0_2320 : std_logic_vector(7 downto 0);
    signal IMA100_3320 : std_logic_vector(7 downto 0);
    signal IMA101_3330 : std_logic_vector(7 downto 0);
    signal IMA102_3340 : std_logic_vector(7 downto 0);
    signal IMA103_3350 : std_logic_vector(7 downto 0);
    signal IMA104_3360 : std_logic_vector(7 downto 0);
    signal IMA105_3370 : std_logic_vector(7 downto 0);
    signal IMA106_3380 : std_logic_vector(7 downto 0);
    signal IMA107_3390 : std_logic_vector(7 downto 0);
    signal IMA108_3400 : std_logic_vector(7 downto 0);
    signal IMA109_3410 : std_logic_vector(7 downto 0);
    signal IMA10_2420 : std_logic_vector(7 downto 0);
    signal IMA110_3420 : std_logic_vector(7 downto 0);
    signal IMA111_3430 : std_logic_vector(7 downto 0);
    signal IMA112_3440 : std_logic_vector(7 downto 0);
    signal IMA113_3450 : std_logic_vector(7 downto 0);
    signal IMA114_3460 : std_logic_vector(7 downto 0);
    signal IMA115_3470 : std_logic_vector(7 downto 0);
    signal IMA116_3480 : std_logic_vector(7 downto 0);
    signal IMA117_3490 : std_logic_vector(7 downto 0);
    signal IMA118_3500 : std_logic_vector(7 downto 0);
    signal IMA119_3510 : std_logic_vector(7 downto 0);
    signal IMA11_2430 : std_logic_vector(7 downto 0);
    signal IMA120_3520 : std_logic_vector(7 downto 0);
    signal IMA121_3530 : std_logic_vector(7 downto 0);
    signal IMA122_3540 : std_logic_vector(7 downto 0);
    signal IMA123_3550 : std_logic_vector(7 downto 0);
    signal IMA124_3560 : std_logic_vector(7 downto 0);
    signal IMA125_3570 : std_logic_vector(7 downto 0);
    signal IMA126_3580 : std_logic_vector(7 downto 0);
    signal IMA127_3590 : std_logic_vector(7 downto 0);
    signal IMA12_2440 : std_logic_vector(7 downto 0);
    signal IMA13_2450 : std_logic_vector(7 downto 0);
    signal IMA14_2460 : std_logic_vector(7 downto 0);
    signal IMA15_2470 : std_logic_vector(7 downto 0);
    signal IMA16_2480 : std_logic_vector(7 downto 0);
    signal IMA17_2490 : std_logic_vector(7 downto 0);
    signal IMA18_2500 : std_logic_vector(7 downto 0);
    signal IMA19_2510 : std_logic_vector(7 downto 0);
    signal IMA1_2330 : std_logic_vector(7 downto 0);
    signal IMA20_2520 : std_logic_vector(7 downto 0);
    signal IMA21_2530 : std_logic_vector(7 downto 0);
    signal IMA22_2540 : std_logic_vector(7 downto 0);
    signal IMA23_2550 : std_logic_vector(7 downto 0);
    signal IMA24_2560 : std_logic_vector(7 downto 0);
    signal IMA25_2570 : std_logic_vector(7 downto 0);
    signal IMA26_2580 : std_logic_vector(7 downto 0);
    signal IMA27_2590 : std_logic_vector(7 downto 0);
    signal IMA28_2600 : std_logic_vector(7 downto 0);
    signal IMA29_2610 : std_logic_vector(7 downto 0);
    signal IMA2_2340 : std_logic_vector(7 downto 0);
    signal IMA30_2620 : std_logic_vector(7 downto 0);
    signal IMA31_2630 : std_logic_vector(7 downto 0);
    signal IMA32_2640 : std_logic_vector(7 downto 0);
    signal IMA33_2650 : std_logic_vector(7 downto 0);
    signal IMA34_2660 : std_logic_vector(7 downto 0);
    signal IMA35_2670 : std_logic_vector(7 downto 0);
    signal IMA36_2680 : std_logic_vector(7 downto 0);
    signal IMA37_2690 : std_logic_vector(7 downto 0);
    signal IMA38_2700 : std_logic_vector(7 downto 0);
    signal IMA39_2710 : std_logic_vector(7 downto 0);
    signal IMA3_2350 : std_logic_vector(7 downto 0);
    signal IMA40_2720 : std_logic_vector(7 downto 0);
    signal IMA41_2730 : std_logic_vector(7 downto 0);
    signal IMA42_2740 : std_logic_vector(7 downto 0);
    signal IMA43_2750 : std_logic_vector(7 downto 0);
    signal IMA44_2760 : std_logic_vector(7 downto 0);
    signal IMA45_2770 : std_logic_vector(7 downto 0);
    signal IMA46_2780 : std_logic_vector(7 downto 0);
    signal IMA47_2790 : std_logic_vector(7 downto 0);
    signal IMA48_2800 : std_logic_vector(7 downto 0);
    signal IMA49_2810 : std_logic_vector(7 downto 0);
    signal IMA4_2360 : std_logic_vector(7 downto 0);
    signal IMA50_2820 : std_logic_vector(7 downto 0);
    signal IMA51_2830 : std_logic_vector(7 downto 0);
    signal IMA52_2840 : std_logic_vector(7 downto 0);
    signal IMA53_2850 : std_logic_vector(7 downto 0);
    signal IMA54_2860 : std_logic_vector(7 downto 0);
    signal IMA55_2870 : std_logic_vector(7 downto 0);
    signal IMA56_2880 : std_logic_vector(7 downto 0);
    signal IMA57_2890 : std_logic_vector(7 downto 0);
    signal IMA58_2900 : std_logic_vector(7 downto 0);
    signal IMA59_2910 : std_logic_vector(7 downto 0);
    signal IMA5_2370 : std_logic_vector(7 downto 0);
    signal IMA60_2920 : std_logic_vector(7 downto 0);
    signal IMA61_2930 : std_logic_vector(7 downto 0);
    signal IMA62_2940 : std_logic_vector(7 downto 0);
    signal IMA63_2950 : std_logic_vector(7 downto 0);
    signal IMA64_2960 : std_logic_vector(7 downto 0);
    signal IMA65_2970 : std_logic_vector(7 downto 0);
    signal IMA66_2980 : std_logic_vector(7 downto 0);
    signal IMA67_2990 : std_logic_vector(7 downto 0);
    signal IMA68_3000 : std_logic_vector(7 downto 0);
    signal IMA69_3010 : std_logic_vector(7 downto 0);
    signal IMA6_2380 : std_logic_vector(7 downto 0);
    signal IMA70_3020 : std_logic_vector(7 downto 0);
    signal IMA71_3030 : std_logic_vector(7 downto 0);
    signal IMA72_3040 : std_logic_vector(7 downto 0);
    signal IMA73_3050 : std_logic_vector(7 downto 0);
    signal IMA74_3060 : std_logic_vector(7 downto 0);
    signal IMA75_3070 : std_logic_vector(7 downto 0);
    signal IMA76_3080 : std_logic_vector(7 downto 0);
    signal IMA77_3090 : std_logic_vector(7 downto 0);
    signal IMA78_3100 : std_logic_vector(7 downto 0);
    signal IMA79_3110 : std_logic_vector(7 downto 0);
    signal IMA7_2390 : std_logic_vector(7 downto 0);
    signal IMA80_3120 : std_logic_vector(7 downto 0);
    signal IMA81_3130 : std_logic_vector(7 downto 0);
    signal IMA82_3140 : std_logic_vector(7 downto 0);
    signal IMA83_3150 : std_logic_vector(7 downto 0);
    signal IMA84_3160 : std_logic_vector(7 downto 0);
    signal IMA85_3170 : std_logic_vector(7 downto 0);
    signal IMA86_3180 : std_logic_vector(7 downto 0);
    signal IMA87_3190 : std_logic_vector(7 downto 0);
    signal IMA88_3200 : std_logic_vector(7 downto 0);
    signal IMA89_3210 : std_logic_vector(7 downto 0);
    signal IMA8_2400 : std_logic_vector(7 downto 0);
    signal IMA90_3220 : std_logic_vector(7 downto 0);
    signal IMA91_3230 : std_logic_vector(7 downto 0);
    signal IMA92_3240 : std_logic_vector(7 downto 0);
    signal IMA93_3250 : std_logic_vector(7 downto 0);
    signal IMA94_3260 : std_logic_vector(7 downto 0);
    signal IMA95_3270 : std_logic_vector(7 downto 0);
    signal IMA96_3280 : std_logic_vector(7 downto 0);
    signal IMA97_3290 : std_logic_vector(7 downto 0);
    signal IMA98_3300 : std_logic_vector(7 downto 0);
    signal IMA99_3310 : std_logic_vector(7 downto 0);
    signal IMA9_2410 : std_logic_vector(7 downto 0);
    signal IMB0_3598 : std_logic_vector(7 downto 0);
    signal IMB10_3678 : std_logic_vector(7 downto 0);
    signal IMB11_3686 : std_logic_vector(7 downto 0);
    signal IMB12_3694 : std_logic_vector(7 downto 0);
    signal IMB13_3702 : std_logic_vector(7 downto 0);
    signal IMB14_3710 : std_logic_vector(7 downto 0);
    signal IMB15_3718 : std_logic_vector(7 downto 0);
    signal IMB16_3726 : std_logic_vector(7 downto 0);
    signal IMB17_3734 : std_logic_vector(7 downto 0);
    signal IMB18_3742 : std_logic_vector(7 downto 0);
    signal IMB19_3750 : std_logic_vector(7 downto 0);
    signal IMB1_3606 : std_logic_vector(7 downto 0);
    signal IMB20_3758 : std_logic_vector(7 downto 0);
    signal IMB21_3766 : std_logic_vector(7 downto 0);
    signal IMB22_3774 : std_logic_vector(7 downto 0);
    signal IMB23_3782 : std_logic_vector(7 downto 0);
    signal IMB24_3790 : std_logic_vector(7 downto 0);
    signal IMB25_3798 : std_logic_vector(7 downto 0);
    signal IMB26_3806 : std_logic_vector(7 downto 0);
    signal IMB27_3814 : std_logic_vector(7 downto 0);
    signal IMB28_3822 : std_logic_vector(7 downto 0);
    signal IMB29_3830 : std_logic_vector(7 downto 0);
    signal IMB2_3614 : std_logic_vector(7 downto 0);
    signal IMB30_3838 : std_logic_vector(7 downto 0);
    signal IMB31_3846 : std_logic_vector(7 downto 0);
    signal IMB32_3854 : std_logic_vector(7 downto 0);
    signal IMB33_3862 : std_logic_vector(7 downto 0);
    signal IMB34_3870 : std_logic_vector(7 downto 0);
    signal IMB35_3878 : std_logic_vector(7 downto 0);
    signal IMB36_3886 : std_logic_vector(7 downto 0);
    signal IMB37_3894 : std_logic_vector(7 downto 0);
    signal IMB38_3902 : std_logic_vector(7 downto 0);
    signal IMB39_3910 : std_logic_vector(7 downto 0);
    signal IMB3_3622 : std_logic_vector(7 downto 0);
    signal IMB40_3918 : std_logic_vector(7 downto 0);
    signal IMB41_3926 : std_logic_vector(7 downto 0);
    signal IMB42_3934 : std_logic_vector(7 downto 0);
    signal IMB43_3942 : std_logic_vector(7 downto 0);
    signal IMB44_3950 : std_logic_vector(7 downto 0);
    signal IMB45_3958 : std_logic_vector(7 downto 0);
    signal IMB46_3966 : std_logic_vector(7 downto 0);
    signal IMB47_3974 : std_logic_vector(7 downto 0);
    signal IMB48_3982 : std_logic_vector(7 downto 0);
    signal IMB49_3990 : std_logic_vector(7 downto 0);
    signal IMB4_3630 : std_logic_vector(7 downto 0);
    signal IMB50_3998 : std_logic_vector(7 downto 0);
    signal IMB51_4006 : std_logic_vector(7 downto 0);
    signal IMB52_4014 : std_logic_vector(7 downto 0);
    signal IMB53_4022 : std_logic_vector(7 downto 0);
    signal IMB54_4030 : std_logic_vector(7 downto 0);
    signal IMB55_4038 : std_logic_vector(7 downto 0);
    signal IMB56_4046 : std_logic_vector(7 downto 0);
    signal IMB57_4054 : std_logic_vector(7 downto 0);
    signal IMB58_4062 : std_logic_vector(7 downto 0);
    signal IMB59_4070 : std_logic_vector(7 downto 0);
    signal IMB5_3638 : std_logic_vector(7 downto 0);
    signal IMB60_4078 : std_logic_vector(7 downto 0);
    signal IMB61_4086 : std_logic_vector(7 downto 0);
    signal IMB62_4094 : std_logic_vector(7 downto 0);
    signal IMB63_4102 : std_logic_vector(7 downto 0);
    signal IMB6_3646 : std_logic_vector(7 downto 0);
    signal IMB7_3654 : std_logic_vector(7 downto 0);
    signal IMB8_3662 : std_logic_vector(7 downto 0);
    signal IMB9_3670 : std_logic_vector(7 downto 0);
    signal IMC0_4110 : std_logic_vector(7 downto 0);
    signal IMC10_4190 : std_logic_vector(7 downto 0);
    signal IMC11_4198 : std_logic_vector(7 downto 0);
    signal IMC12_4206 : std_logic_vector(7 downto 0);
    signal IMC13_4214 : std_logic_vector(7 downto 0);
    signal IMC14_4222 : std_logic_vector(7 downto 0);
    signal IMC15_4230 : std_logic_vector(7 downto 0);
    signal IMC16_4238 : std_logic_vector(7 downto 0);
    signal IMC17_4246 : std_logic_vector(7 downto 0);
    signal IMC18_4254 : std_logic_vector(7 downto 0);
    signal IMC19_4262 : std_logic_vector(7 downto 0);
    signal IMC1_4118 : std_logic_vector(7 downto 0);
    signal IMC20_4270 : std_logic_vector(7 downto 0);
    signal IMC21_4278 : std_logic_vector(7 downto 0);
    signal IMC22_4286 : std_logic_vector(7 downto 0);
    signal IMC23_4294 : std_logic_vector(7 downto 0);
    signal IMC24_4302 : std_logic_vector(7 downto 0);
    signal IMC25_4310 : std_logic_vector(7 downto 0);
    signal IMC26_4318 : std_logic_vector(7 downto 0);
    signal IMC27_4326 : std_logic_vector(7 downto 0);
    signal IMC28_4334 : std_logic_vector(7 downto 0);
    signal IMC29_4342 : std_logic_vector(7 downto 0);
    signal IMC2_4126 : std_logic_vector(7 downto 0);
    signal IMC30_4350 : std_logic_vector(7 downto 0);
    signal IMC31_4358 : std_logic_vector(7 downto 0);
    signal IMC3_4134 : std_logic_vector(7 downto 0);
    signal IMC4_4142 : std_logic_vector(7 downto 0);
    signal IMC5_4150 : std_logic_vector(7 downto 0);
    signal IMC6_4158 : std_logic_vector(7 downto 0);
    signal IMC7_4166 : std_logic_vector(7 downto 0);
    signal IMC8_4174 : std_logic_vector(7 downto 0);
    signal IMC9_4182 : std_logic_vector(7 downto 0);
    signal IMD0_4366 : std_logic_vector(7 downto 0);
    signal IMD10_4446 : std_logic_vector(7 downto 0);
    signal IMD11_4454 : std_logic_vector(7 downto 0);
    signal IMD12_4462 : std_logic_vector(7 downto 0);
    signal IMD13_4470 : std_logic_vector(7 downto 0);
    signal IMD14_4478 : std_logic_vector(7 downto 0);
    signal IMD15_4486 : std_logic_vector(7 downto 0);
    signal IMD1_4374 : std_logic_vector(7 downto 0);
    signal IMD2_4382 : std_logic_vector(7 downto 0);
    signal IMD3_4390 : std_logic_vector(7 downto 0);
    signal IMD4_4398 : std_logic_vector(7 downto 0);
    signal IMD5_4406 : std_logic_vector(7 downto 0);
    signal IMD6_4414 : std_logic_vector(7 downto 0);
    signal IMD7_4422 : std_logic_vector(7 downto 0);
    signal IMD8_4430 : std_logic_vector(7 downto 0);
    signal IMD9_4438 : std_logic_vector(7 downto 0);
    signal IME0_4494 : std_logic_vector(7 downto 0);
    signal IME1_4502 : std_logic_vector(7 downto 0);
    signal IME2_4510 : std_logic_vector(7 downto 0);
    signal IME3_4518 : std_logic_vector(7 downto 0);
    signal IME4_4526 : std_logic_vector(7 downto 0);
    signal IME5_4534 : std_logic_vector(7 downto 0);
    signal IME6_4542 : std_logic_vector(7 downto 0);
    signal IME7_4550 : std_logic_vector(7 downto 0);
    signal IMF0_4558 : std_logic_vector(7 downto 0);
    signal IMF1_4566 : std_logic_vector(7 downto 0);
    signal IMF2_4574 : std_logic_vector(7 downto 0);
    signal IMF3_4582 : std_logic_vector(7 downto 0);
    signal IMG0_4590 : std_logic_vector(7 downto 0);
    signal IMG1_4598 : std_logic_vector(7 downto 0);
    signal konst_2313_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2323_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2333_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2343_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2353_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2363_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2373_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2383_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2393_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2403_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2413_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2423_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2433_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2443_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2453_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2463_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2473_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2483_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2493_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2503_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2513_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2523_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2533_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2543_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2553_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2563_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2573_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2583_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2593_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2603_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2613_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2623_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2633_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2643_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2653_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2663_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2673_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2683_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2693_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2703_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2713_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2723_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2733_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2743_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2753_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2763_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2773_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2783_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2793_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2803_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2813_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2823_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2833_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2843_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2853_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2863_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2873_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2883_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2893_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2903_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2913_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2923_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2933_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2943_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2953_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2963_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2973_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2983_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2993_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3003_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3013_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3023_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3033_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3043_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3053_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3063_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3073_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3083_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3093_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3103_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3113_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3123_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3133_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3143_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3153_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3163_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3173_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3183_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3193_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3203_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3213_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3223_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3233_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3243_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3253_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3263_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3273_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3283_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3293_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3303_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3313_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3323_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3333_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3343_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3353_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3363_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3373_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3383_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3393_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3403_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3413_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3423_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3433_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3443_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3453_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3463_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3473_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3483_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3493_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3503_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3513_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3523_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3533_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3543_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3553_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3563_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3573_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3583_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3593_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3601_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3609_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3617_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3625_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3633_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3641_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3649_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3657_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3665_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3673_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3681_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3689_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3697_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3705_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3713_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3721_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3729_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3737_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3745_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3753_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3761_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3769_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3777_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3785_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3793_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3801_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3809_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3817_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3825_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3833_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3841_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3849_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3857_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3865_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3873_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3881_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3889_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3897_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3905_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3913_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3921_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3929_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3937_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3945_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3953_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3961_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3969_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3977_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3985_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3993_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4001_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4009_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4017_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4025_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4033_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4041_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4049_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4057_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4065_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4073_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4081_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4089_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4097_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4105_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4113_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4121_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4129_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4137_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4145_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4153_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4161_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4169_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4177_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4185_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4193_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4201_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4209_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4217_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4225_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4233_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4241_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4249_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4257_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4265_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4273_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4281_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4289_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4297_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4305_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4313_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4321_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4329_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4337_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4345_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4353_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4361_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4369_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4377_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4385_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4393_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4401_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4409_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4417_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4425_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4433_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4441_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4449_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4457_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4465_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4473_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4481_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4489_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4497_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4505_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4513_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4521_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4529_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4537_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4545_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4553_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4561_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4569_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4577_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4585_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4593_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4601_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2316_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2318_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2326_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2328_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2336_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2338_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2346_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2348_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2356_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2358_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2366_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2368_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2376_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2378_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2386_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2388_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2396_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2398_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2406_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2408_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2416_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2418_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2426_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2428_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2436_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2438_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2446_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2448_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2456_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2458_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2466_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2468_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2476_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2478_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2486_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2488_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2496_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2498_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2506_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2508_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2516_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2518_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2526_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2528_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2536_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2538_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2546_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2548_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2556_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2558_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2566_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2568_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2576_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2578_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2586_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2588_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2596_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2598_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2606_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2608_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2616_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2618_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2626_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2628_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2636_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2638_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2646_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2648_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2656_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2658_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2666_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2668_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2676_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2678_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2686_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2688_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2696_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2698_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2706_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2708_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2716_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2718_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2726_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2728_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2736_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2738_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2746_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2748_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2756_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2758_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2766_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2768_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2776_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2778_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2786_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2788_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2796_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2798_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2806_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2808_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2816_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2818_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2826_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2828_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2836_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2838_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2846_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2848_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2856_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2858_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2866_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2868_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2876_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2878_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2886_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2888_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2896_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2898_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2906_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2908_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2916_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2918_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2926_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2928_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2936_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2938_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2946_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2948_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2956_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2958_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2966_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2968_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2976_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2978_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2986_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2988_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2996_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2998_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3006_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3008_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3016_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3018_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3026_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3028_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3036_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3038_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3046_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3048_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3056_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3058_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3066_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3068_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3076_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3078_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3086_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3088_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3096_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3098_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3106_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3108_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3116_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3118_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3126_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3128_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3136_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3138_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3146_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3148_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3156_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3158_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3166_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3168_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3176_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3178_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3186_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3188_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3196_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3198_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3206_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3208_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3216_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3218_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3226_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3228_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3236_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3238_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3246_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3248_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3256_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3258_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3266_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3268_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3276_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3278_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3286_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3288_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3296_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3298_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3306_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3308_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3316_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3318_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3326_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3328_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3336_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3338_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3346_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3348_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3356_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3358_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3366_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3368_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3376_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3378_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3386_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3388_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3396_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3398_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3406_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3408_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3416_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3418_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3426_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3428_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3436_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3438_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3446_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3448_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3456_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3458_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3466_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3468_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3476_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3478_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3486_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3488_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3496_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3498_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3506_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3508_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3516_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3518_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3526_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3528_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3536_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3538_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3546_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3548_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3556_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3558_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3566_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3568_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3576_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3578_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3586_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3588_wire_constant : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    konst_2313_wire_constant <= "00000000";
    konst_2323_wire_constant <= "00000000";
    konst_2333_wire_constant <= "00000000";
    konst_2343_wire_constant <= "00000000";
    konst_2353_wire_constant <= "00000000";
    konst_2363_wire_constant <= "00000000";
    konst_2373_wire_constant <= "00000000";
    konst_2383_wire_constant <= "00000000";
    konst_2393_wire_constant <= "00000000";
    konst_2403_wire_constant <= "00000000";
    konst_2413_wire_constant <= "00000000";
    konst_2423_wire_constant <= "00000000";
    konst_2433_wire_constant <= "00000000";
    konst_2443_wire_constant <= "00000000";
    konst_2453_wire_constant <= "00000000";
    konst_2463_wire_constant <= "00000000";
    konst_2473_wire_constant <= "00000000";
    konst_2483_wire_constant <= "00000000";
    konst_2493_wire_constant <= "00000000";
    konst_2503_wire_constant <= "00000000";
    konst_2513_wire_constant <= "00000000";
    konst_2523_wire_constant <= "00000000";
    konst_2533_wire_constant <= "00000000";
    konst_2543_wire_constant <= "00000000";
    konst_2553_wire_constant <= "00000000";
    konst_2563_wire_constant <= "00000000";
    konst_2573_wire_constant <= "00000000";
    konst_2583_wire_constant <= "00000000";
    konst_2593_wire_constant <= "00000000";
    konst_2603_wire_constant <= "00000000";
    konst_2613_wire_constant <= "00000000";
    konst_2623_wire_constant <= "00000000";
    konst_2633_wire_constant <= "00000000";
    konst_2643_wire_constant <= "00000000";
    konst_2653_wire_constant <= "00000000";
    konst_2663_wire_constant <= "00000000";
    konst_2673_wire_constant <= "00000000";
    konst_2683_wire_constant <= "00000000";
    konst_2693_wire_constant <= "00000000";
    konst_2703_wire_constant <= "00000000";
    konst_2713_wire_constant <= "00000000";
    konst_2723_wire_constant <= "00000000";
    konst_2733_wire_constant <= "00000000";
    konst_2743_wire_constant <= "00000000";
    konst_2753_wire_constant <= "00000000";
    konst_2763_wire_constant <= "00000000";
    konst_2773_wire_constant <= "00000000";
    konst_2783_wire_constant <= "00000000";
    konst_2793_wire_constant <= "00000000";
    konst_2803_wire_constant <= "00000000";
    konst_2813_wire_constant <= "00000000";
    konst_2823_wire_constant <= "00000000";
    konst_2833_wire_constant <= "00000000";
    konst_2843_wire_constant <= "00000000";
    konst_2853_wire_constant <= "00000000";
    konst_2863_wire_constant <= "00000000";
    konst_2873_wire_constant <= "00000000";
    konst_2883_wire_constant <= "00000000";
    konst_2893_wire_constant <= "00000000";
    konst_2903_wire_constant <= "00000000";
    konst_2913_wire_constant <= "00000000";
    konst_2923_wire_constant <= "00000000";
    konst_2933_wire_constant <= "00000000";
    konst_2943_wire_constant <= "00000000";
    konst_2953_wire_constant <= "00000000";
    konst_2963_wire_constant <= "00000000";
    konst_2973_wire_constant <= "00000000";
    konst_2983_wire_constant <= "00000000";
    konst_2993_wire_constant <= "00000000";
    konst_3003_wire_constant <= "00000000";
    konst_3013_wire_constant <= "00000000";
    konst_3023_wire_constant <= "00000000";
    konst_3033_wire_constant <= "00000000";
    konst_3043_wire_constant <= "00000000";
    konst_3053_wire_constant <= "00000000";
    konst_3063_wire_constant <= "00000000";
    konst_3073_wire_constant <= "00000000";
    konst_3083_wire_constant <= "00000000";
    konst_3093_wire_constant <= "00000000";
    konst_3103_wire_constant <= "00000000";
    konst_3113_wire_constant <= "00000000";
    konst_3123_wire_constant <= "00000000";
    konst_3133_wire_constant <= "00000000";
    konst_3143_wire_constant <= "00000000";
    konst_3153_wire_constant <= "00000000";
    konst_3163_wire_constant <= "00000000";
    konst_3173_wire_constant <= "00000000";
    konst_3183_wire_constant <= "00000000";
    konst_3193_wire_constant <= "00000000";
    konst_3203_wire_constant <= "00000000";
    konst_3213_wire_constant <= "00000000";
    konst_3223_wire_constant <= "00000000";
    konst_3233_wire_constant <= "00000000";
    konst_3243_wire_constant <= "00000000";
    konst_3253_wire_constant <= "00000000";
    konst_3263_wire_constant <= "00000000";
    konst_3273_wire_constant <= "00000000";
    konst_3283_wire_constant <= "00000000";
    konst_3293_wire_constant <= "00000000";
    konst_3303_wire_constant <= "00000000";
    konst_3313_wire_constant <= "00000000";
    konst_3323_wire_constant <= "00000000";
    konst_3333_wire_constant <= "00000000";
    konst_3343_wire_constant <= "00000000";
    konst_3353_wire_constant <= "00000000";
    konst_3363_wire_constant <= "00000000";
    konst_3373_wire_constant <= "00000000";
    konst_3383_wire_constant <= "00000000";
    konst_3393_wire_constant <= "00000000";
    konst_3403_wire_constant <= "00000000";
    konst_3413_wire_constant <= "00000000";
    konst_3423_wire_constant <= "00000000";
    konst_3433_wire_constant <= "00000000";
    konst_3443_wire_constant <= "00000000";
    konst_3453_wire_constant <= "00000000";
    konst_3463_wire_constant <= "00000000";
    konst_3473_wire_constant <= "00000000";
    konst_3483_wire_constant <= "00000000";
    konst_3493_wire_constant <= "00000000";
    konst_3503_wire_constant <= "00000000";
    konst_3513_wire_constant <= "00000000";
    konst_3523_wire_constant <= "00000000";
    konst_3533_wire_constant <= "00000000";
    konst_3543_wire_constant <= "00000000";
    konst_3553_wire_constant <= "00000000";
    konst_3563_wire_constant <= "00000000";
    konst_3573_wire_constant <= "00000000";
    konst_3583_wire_constant <= "00000000";
    konst_3593_wire_constant <= "00000001";
    konst_3601_wire_constant <= "00000001";
    konst_3609_wire_constant <= "00000001";
    konst_3617_wire_constant <= "00000001";
    konst_3625_wire_constant <= "00000001";
    konst_3633_wire_constant <= "00000001";
    konst_3641_wire_constant <= "00000001";
    konst_3649_wire_constant <= "00000001";
    konst_3657_wire_constant <= "00000001";
    konst_3665_wire_constant <= "00000001";
    konst_3673_wire_constant <= "00000001";
    konst_3681_wire_constant <= "00000001";
    konst_3689_wire_constant <= "00000001";
    konst_3697_wire_constant <= "00000001";
    konst_3705_wire_constant <= "00000001";
    konst_3713_wire_constant <= "00000001";
    konst_3721_wire_constant <= "00000001";
    konst_3729_wire_constant <= "00000001";
    konst_3737_wire_constant <= "00000001";
    konst_3745_wire_constant <= "00000001";
    konst_3753_wire_constant <= "00000001";
    konst_3761_wire_constant <= "00000001";
    konst_3769_wire_constant <= "00000001";
    konst_3777_wire_constant <= "00000001";
    konst_3785_wire_constant <= "00000001";
    konst_3793_wire_constant <= "00000001";
    konst_3801_wire_constant <= "00000001";
    konst_3809_wire_constant <= "00000001";
    konst_3817_wire_constant <= "00000001";
    konst_3825_wire_constant <= "00000001";
    konst_3833_wire_constant <= "00000001";
    konst_3841_wire_constant <= "00000001";
    konst_3849_wire_constant <= "00000001";
    konst_3857_wire_constant <= "00000001";
    konst_3865_wire_constant <= "00000001";
    konst_3873_wire_constant <= "00000001";
    konst_3881_wire_constant <= "00000001";
    konst_3889_wire_constant <= "00000001";
    konst_3897_wire_constant <= "00000001";
    konst_3905_wire_constant <= "00000001";
    konst_3913_wire_constant <= "00000001";
    konst_3921_wire_constant <= "00000001";
    konst_3929_wire_constant <= "00000001";
    konst_3937_wire_constant <= "00000001";
    konst_3945_wire_constant <= "00000001";
    konst_3953_wire_constant <= "00000001";
    konst_3961_wire_constant <= "00000001";
    konst_3969_wire_constant <= "00000001";
    konst_3977_wire_constant <= "00000001";
    konst_3985_wire_constant <= "00000001";
    konst_3993_wire_constant <= "00000001";
    konst_4001_wire_constant <= "00000001";
    konst_4009_wire_constant <= "00000001";
    konst_4017_wire_constant <= "00000001";
    konst_4025_wire_constant <= "00000001";
    konst_4033_wire_constant <= "00000001";
    konst_4041_wire_constant <= "00000001";
    konst_4049_wire_constant <= "00000001";
    konst_4057_wire_constant <= "00000001";
    konst_4065_wire_constant <= "00000001";
    konst_4073_wire_constant <= "00000001";
    konst_4081_wire_constant <= "00000001";
    konst_4089_wire_constant <= "00000001";
    konst_4097_wire_constant <= "00000001";
    konst_4105_wire_constant <= "00000010";
    konst_4113_wire_constant <= "00000010";
    konst_4121_wire_constant <= "00000010";
    konst_4129_wire_constant <= "00000010";
    konst_4137_wire_constant <= "00000010";
    konst_4145_wire_constant <= "00000010";
    konst_4153_wire_constant <= "00000010";
    konst_4161_wire_constant <= "00000010";
    konst_4169_wire_constant <= "00000010";
    konst_4177_wire_constant <= "00000010";
    konst_4185_wire_constant <= "00000010";
    konst_4193_wire_constant <= "00000010";
    konst_4201_wire_constant <= "00000010";
    konst_4209_wire_constant <= "00000010";
    konst_4217_wire_constant <= "00000010";
    konst_4225_wire_constant <= "00000010";
    konst_4233_wire_constant <= "00000010";
    konst_4241_wire_constant <= "00000010";
    konst_4249_wire_constant <= "00000010";
    konst_4257_wire_constant <= "00000010";
    konst_4265_wire_constant <= "00000010";
    konst_4273_wire_constant <= "00000010";
    konst_4281_wire_constant <= "00000010";
    konst_4289_wire_constant <= "00000010";
    konst_4297_wire_constant <= "00000010";
    konst_4305_wire_constant <= "00000010";
    konst_4313_wire_constant <= "00000010";
    konst_4321_wire_constant <= "00000010";
    konst_4329_wire_constant <= "00000010";
    konst_4337_wire_constant <= "00000010";
    konst_4345_wire_constant <= "00000010";
    konst_4353_wire_constant <= "00000010";
    konst_4361_wire_constant <= "00000011";
    konst_4369_wire_constant <= "00000011";
    konst_4377_wire_constant <= "00000011";
    konst_4385_wire_constant <= "00000011";
    konst_4393_wire_constant <= "00000011";
    konst_4401_wire_constant <= "00000011";
    konst_4409_wire_constant <= "00000011";
    konst_4417_wire_constant <= "00000011";
    konst_4425_wire_constant <= "00000011";
    konst_4433_wire_constant <= "00000011";
    konst_4441_wire_constant <= "00000011";
    konst_4449_wire_constant <= "00000011";
    konst_4457_wire_constant <= "00000011";
    konst_4465_wire_constant <= "00000011";
    konst_4473_wire_constant <= "00000011";
    konst_4481_wire_constant <= "00000011";
    konst_4489_wire_constant <= "00000100";
    konst_4497_wire_constant <= "00000100";
    konst_4505_wire_constant <= "00000100";
    konst_4513_wire_constant <= "00000100";
    konst_4521_wire_constant <= "00000100";
    konst_4529_wire_constant <= "00000100";
    konst_4537_wire_constant <= "00000100";
    konst_4545_wire_constant <= "00000100";
    konst_4553_wire_constant <= "00000101";
    konst_4561_wire_constant <= "00000101";
    konst_4569_wire_constant <= "00000101";
    konst_4577_wire_constant <= "00000101";
    konst_4585_wire_constant <= "00000110";
    konst_4593_wire_constant <= "00000110";
    konst_4601_wire_constant <= "00000111";
    type_cast_2316_wire_constant <= "00001001";
    type_cast_2318_wire_constant <= "01010010";
    type_cast_2326_wire_constant <= "11010101";
    type_cast_2328_wire_constant <= "01101010";
    type_cast_2336_wire_constant <= "00110110";
    type_cast_2338_wire_constant <= "00110000";
    type_cast_2346_wire_constant <= "00111000";
    type_cast_2348_wire_constant <= "10100101";
    type_cast_2356_wire_constant <= "01000000";
    type_cast_2358_wire_constant <= "10111111";
    type_cast_2366_wire_constant <= "10011110";
    type_cast_2368_wire_constant <= "10100011";
    type_cast_2376_wire_constant <= "11110011";
    type_cast_2378_wire_constant <= "10000001";
    type_cast_2386_wire_constant <= "11111011";
    type_cast_2388_wire_constant <= "11010111";
    type_cast_2396_wire_constant <= "11100011";
    type_cast_2398_wire_constant <= "01111100";
    type_cast_2406_wire_constant <= "10000010";
    type_cast_2408_wire_constant <= "00111001";
    type_cast_2416_wire_constant <= "00101111";
    type_cast_2418_wire_constant <= "10011011";
    type_cast_2426_wire_constant <= "10000111";
    type_cast_2428_wire_constant <= "11111111";
    type_cast_2436_wire_constant <= "10001110";
    type_cast_2438_wire_constant <= "00110100";
    type_cast_2446_wire_constant <= "01000100";
    type_cast_2448_wire_constant <= "01000011";
    type_cast_2456_wire_constant <= "11011110";
    type_cast_2458_wire_constant <= "11000100";
    type_cast_2466_wire_constant <= "11001011";
    type_cast_2468_wire_constant <= "11101001";
    type_cast_2476_wire_constant <= "01111011";
    type_cast_2478_wire_constant <= "01010100";
    type_cast_2486_wire_constant <= "00110010";
    type_cast_2488_wire_constant <= "10010100";
    type_cast_2496_wire_constant <= "11000010";
    type_cast_2498_wire_constant <= "10100110";
    type_cast_2506_wire_constant <= "00111101";
    type_cast_2508_wire_constant <= "00100011";
    type_cast_2516_wire_constant <= "01001100";
    type_cast_2518_wire_constant <= "11101110";
    type_cast_2526_wire_constant <= "00001011";
    type_cast_2528_wire_constant <= "10010101";
    type_cast_2536_wire_constant <= "11111010";
    type_cast_2538_wire_constant <= "01000010";
    type_cast_2546_wire_constant <= "01001110";
    type_cast_2548_wire_constant <= "11000011";
    type_cast_2556_wire_constant <= "00101110";
    type_cast_2558_wire_constant <= "00001000";
    type_cast_2566_wire_constant <= "01100110";
    type_cast_2568_wire_constant <= "10100001";
    type_cast_2576_wire_constant <= "11011001";
    type_cast_2578_wire_constant <= "00101000";
    type_cast_2586_wire_constant <= "10110010";
    type_cast_2588_wire_constant <= "00100100";
    type_cast_2596_wire_constant <= "01011011";
    type_cast_2598_wire_constant <= "01110110";
    type_cast_2606_wire_constant <= "01001001";
    type_cast_2608_wire_constant <= "10100010";
    type_cast_2616_wire_constant <= "10001011";
    type_cast_2618_wire_constant <= "01101101";
    type_cast_2626_wire_constant <= "00100101";
    type_cast_2628_wire_constant <= "11010001";
    type_cast_2636_wire_constant <= "11111000";
    type_cast_2638_wire_constant <= "01110010";
    type_cast_2646_wire_constant <= "01100100";
    type_cast_2648_wire_constant <= "11110110";
    type_cast_2656_wire_constant <= "01101000";
    type_cast_2658_wire_constant <= "10000110";
    type_cast_2666_wire_constant <= "00010110";
    type_cast_2668_wire_constant <= "10011000";
    type_cast_2676_wire_constant <= "10100100";
    type_cast_2678_wire_constant <= "11010100";
    type_cast_2686_wire_constant <= "11001100";
    type_cast_2688_wire_constant <= "01011100";
    type_cast_2696_wire_constant <= "01100101";
    type_cast_2698_wire_constant <= "01011101";
    type_cast_2706_wire_constant <= "10010010";
    type_cast_2708_wire_constant <= "10110110";
    type_cast_2716_wire_constant <= "01110000";
    type_cast_2718_wire_constant <= "01101100";
    type_cast_2726_wire_constant <= "01010000";
    type_cast_2728_wire_constant <= "01001000";
    type_cast_2736_wire_constant <= "11101101";
    type_cast_2738_wire_constant <= "11111101";
    type_cast_2746_wire_constant <= "11011010";
    type_cast_2748_wire_constant <= "10111001";
    type_cast_2756_wire_constant <= "00010101";
    type_cast_2758_wire_constant <= "01011110";
    type_cast_2766_wire_constant <= "01010111";
    type_cast_2768_wire_constant <= "01000110";
    type_cast_2776_wire_constant <= "10001101";
    type_cast_2778_wire_constant <= "10100111";
    type_cast_2786_wire_constant <= "10000100";
    type_cast_2788_wire_constant <= "10011101";
    type_cast_2796_wire_constant <= "11011000";
    type_cast_2798_wire_constant <= "10010000";
    type_cast_2806_wire_constant <= "00000000";
    type_cast_2808_wire_constant <= "10101011";
    type_cast_2816_wire_constant <= "10111100";
    type_cast_2818_wire_constant <= "10001100";
    type_cast_2826_wire_constant <= "00001010";
    type_cast_2828_wire_constant <= "11010011";
    type_cast_2836_wire_constant <= "11100100";
    type_cast_2838_wire_constant <= "11110111";
    type_cast_2846_wire_constant <= "00000101";
    type_cast_2848_wire_constant <= "01011000";
    type_cast_2856_wire_constant <= "10110011";
    type_cast_2858_wire_constant <= "10111000";
    type_cast_2866_wire_constant <= "00000110";
    type_cast_2868_wire_constant <= "01000101";
    type_cast_2876_wire_constant <= "00101100";
    type_cast_2878_wire_constant <= "11010000";
    type_cast_2886_wire_constant <= "10001111";
    type_cast_2888_wire_constant <= "00011110";
    type_cast_2896_wire_constant <= "00111111";
    type_cast_2898_wire_constant <= "11001010";
    type_cast_2906_wire_constant <= "00000010";
    type_cast_2908_wire_constant <= "00001111";
    type_cast_2916_wire_constant <= "10101111";
    type_cast_2918_wire_constant <= "11000001";
    type_cast_2926_wire_constant <= "00000011";
    type_cast_2928_wire_constant <= "10111101";
    type_cast_2936_wire_constant <= "00010011";
    type_cast_2938_wire_constant <= "00000001";
    type_cast_2946_wire_constant <= "01101011";
    type_cast_2948_wire_constant <= "10001010";
    type_cast_2956_wire_constant <= "10010001";
    type_cast_2958_wire_constant <= "00111010";
    type_cast_2966_wire_constant <= "01000001";
    type_cast_2968_wire_constant <= "00010001";
    type_cast_2976_wire_constant <= "01100111";
    type_cast_2978_wire_constant <= "01001111";
    type_cast_2986_wire_constant <= "11101010";
    type_cast_2988_wire_constant <= "11011100";
    type_cast_2996_wire_constant <= "11110010";
    type_cast_2998_wire_constant <= "10010111";
    type_cast_3006_wire_constant <= "11001110";
    type_cast_3008_wire_constant <= "11001111";
    type_cast_3016_wire_constant <= "10110100";
    type_cast_3018_wire_constant <= "11110000";
    type_cast_3026_wire_constant <= "01110011";
    type_cast_3028_wire_constant <= "11100110";
    type_cast_3036_wire_constant <= "10101100";
    type_cast_3038_wire_constant <= "10010110";
    type_cast_3046_wire_constant <= "00100010";
    type_cast_3048_wire_constant <= "01110100";
    type_cast_3056_wire_constant <= "10101101";
    type_cast_3058_wire_constant <= "11100111";
    type_cast_3066_wire_constant <= "10000101";
    type_cast_3068_wire_constant <= "00110101";
    type_cast_3076_wire_constant <= "11111001";
    type_cast_3078_wire_constant <= "11100010";
    type_cast_3086_wire_constant <= "11101000";
    type_cast_3088_wire_constant <= "00110111";
    type_cast_3096_wire_constant <= "01110101";
    type_cast_3098_wire_constant <= "00011100";
    type_cast_3106_wire_constant <= "01101110";
    type_cast_3108_wire_constant <= "11011111";
    type_cast_3116_wire_constant <= "11110001";
    type_cast_3118_wire_constant <= "01000111";
    type_cast_3126_wire_constant <= "01110001";
    type_cast_3128_wire_constant <= "00011010";
    type_cast_3136_wire_constant <= "00101001";
    type_cast_3138_wire_constant <= "00011101";
    type_cast_3146_wire_constant <= "10001001";
    type_cast_3148_wire_constant <= "11000101";
    type_cast_3156_wire_constant <= "10110111";
    type_cast_3158_wire_constant <= "01101111";
    type_cast_3166_wire_constant <= "00001110";
    type_cast_3168_wire_constant <= "01100010";
    type_cast_3176_wire_constant <= "00011000";
    type_cast_3178_wire_constant <= "10101010";
    type_cast_3186_wire_constant <= "00011011";
    type_cast_3188_wire_constant <= "10111110";
    type_cast_3196_wire_constant <= "01010110";
    type_cast_3198_wire_constant <= "11111100";
    type_cast_3206_wire_constant <= "01001011";
    type_cast_3208_wire_constant <= "00111110";
    type_cast_3216_wire_constant <= "11010010";
    type_cast_3218_wire_constant <= "11000110";
    type_cast_3226_wire_constant <= "00100000";
    type_cast_3228_wire_constant <= "01111001";
    type_cast_3236_wire_constant <= "11011011";
    type_cast_3238_wire_constant <= "10011010";
    type_cast_3246_wire_constant <= "11111110";
    type_cast_3248_wire_constant <= "11000000";
    type_cast_3256_wire_constant <= "11001101";
    type_cast_3258_wire_constant <= "01111000";
    type_cast_3266_wire_constant <= "11110100";
    type_cast_3268_wire_constant <= "01011010";
    type_cast_3276_wire_constant <= "11011101";
    type_cast_3278_wire_constant <= "00011111";
    type_cast_3286_wire_constant <= "00110011";
    type_cast_3288_wire_constant <= "10101000";
    type_cast_3296_wire_constant <= "00000111";
    type_cast_3298_wire_constant <= "10001000";
    type_cast_3306_wire_constant <= "00110001";
    type_cast_3308_wire_constant <= "11000111";
    type_cast_3316_wire_constant <= "00010010";
    type_cast_3318_wire_constant <= "10110001";
    type_cast_3326_wire_constant <= "01011001";
    type_cast_3328_wire_constant <= "00010000";
    type_cast_3336_wire_constant <= "10000000";
    type_cast_3338_wire_constant <= "00100111";
    type_cast_3346_wire_constant <= "01011111";
    type_cast_3348_wire_constant <= "11101100";
    type_cast_3356_wire_constant <= "01010001";
    type_cast_3358_wire_constant <= "01100000";
    type_cast_3366_wire_constant <= "10101001";
    type_cast_3368_wire_constant <= "01111111";
    type_cast_3376_wire_constant <= "10110101";
    type_cast_3378_wire_constant <= "00011001";
    type_cast_3386_wire_constant <= "00001101";
    type_cast_3388_wire_constant <= "01001010";
    type_cast_3396_wire_constant <= "11100101";
    type_cast_3398_wire_constant <= "00101101";
    type_cast_3406_wire_constant <= "10011111";
    type_cast_3408_wire_constant <= "01111010";
    type_cast_3416_wire_constant <= "11001001";
    type_cast_3418_wire_constant <= "10010011";
    type_cast_3426_wire_constant <= "11101111";
    type_cast_3428_wire_constant <= "10011100";
    type_cast_3436_wire_constant <= "11100000";
    type_cast_3438_wire_constant <= "10100000";
    type_cast_3446_wire_constant <= "01001101";
    type_cast_3448_wire_constant <= "00111011";
    type_cast_3456_wire_constant <= "00101010";
    type_cast_3458_wire_constant <= "10101110";
    type_cast_3466_wire_constant <= "10110000";
    type_cast_3468_wire_constant <= "11110101";
    type_cast_3476_wire_constant <= "11101011";
    type_cast_3478_wire_constant <= "11001000";
    type_cast_3486_wire_constant <= "00111100";
    type_cast_3488_wire_constant <= "10111011";
    type_cast_3496_wire_constant <= "01010011";
    type_cast_3498_wire_constant <= "10000011";
    type_cast_3506_wire_constant <= "01100001";
    type_cast_3508_wire_constant <= "10011001";
    type_cast_3516_wire_constant <= "00101011";
    type_cast_3518_wire_constant <= "00010111";
    type_cast_3526_wire_constant <= "01111110";
    type_cast_3528_wire_constant <= "00000100";
    type_cast_3536_wire_constant <= "01110111";
    type_cast_3538_wire_constant <= "10111010";
    type_cast_3546_wire_constant <= "00100110";
    type_cast_3548_wire_constant <= "11010110";
    type_cast_3556_wire_constant <= "01101001";
    type_cast_3558_wire_constant <= "11100001";
    type_cast_3566_wire_constant <= "01100011";
    type_cast_3568_wire_constant <= "00010100";
    type_cast_3576_wire_constant <= "00100001";
    type_cast_3578_wire_constant <= "01010101";
    type_cast_3586_wire_constant <= "01111101";
    type_cast_3588_wire_constant <= "00001100";
    -- logger for split-operator MUX_2319_inst flow-through 
    process(IMA0_2320) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_2319_inst:flowthrough inputs: " & " BITSEL_u8_u1_2314_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_2314_wire) & " type_cast_2316_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2316_wire_constant) & " type_cast_2318_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2318_wire_constant) & " outputs:" & " IMA0_2320= "  & Convert_SLV_To_Hex_String(IMA0_2320));
      --
    end process; 
    -- flow-through select operator MUX_2319_inst
    IMA0_2320 <= type_cast_2316_wire_constant when (BITSEL_u8_u1_2314_wire(0) /=  '0') else type_cast_2318_wire_constant;
    -- logger for split-operator MUX_2329_inst flow-through 
    process(IMA1_2330) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_2329_inst:flowthrough inputs: " & " BITSEL_u8_u1_2324_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_2324_wire) & " type_cast_2326_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2326_wire_constant) & " type_cast_2328_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2328_wire_constant) & " outputs:" & " IMA1_2330= "  & Convert_SLV_To_Hex_String(IMA1_2330));
      --
    end process; 
    -- flow-through select operator MUX_2329_inst
    IMA1_2330 <= type_cast_2326_wire_constant when (BITSEL_u8_u1_2324_wire(0) /=  '0') else type_cast_2328_wire_constant;
    -- logger for split-operator MUX_2339_inst flow-through 
    process(IMA2_2340) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_2339_inst:flowthrough inputs: " & " BITSEL_u8_u1_2334_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_2334_wire) & " type_cast_2336_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2336_wire_constant) & " type_cast_2338_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2338_wire_constant) & " outputs:" & " IMA2_2340= "  & Convert_SLV_To_Hex_String(IMA2_2340));
      --
    end process; 
    -- flow-through select operator MUX_2339_inst
    IMA2_2340 <= type_cast_2336_wire_constant when (BITSEL_u8_u1_2334_wire(0) /=  '0') else type_cast_2338_wire_constant;
    -- logger for split-operator MUX_2349_inst flow-through 
    process(IMA3_2350) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_2349_inst:flowthrough inputs: " & " BITSEL_u8_u1_2344_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_2344_wire) & " type_cast_2346_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2346_wire_constant) & " type_cast_2348_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2348_wire_constant) & " outputs:" & " IMA3_2350= "  & Convert_SLV_To_Hex_String(IMA3_2350));
      --
    end process; 
    -- flow-through select operator MUX_2349_inst
    IMA3_2350 <= type_cast_2346_wire_constant when (BITSEL_u8_u1_2344_wire(0) /=  '0') else type_cast_2348_wire_constant;
    -- logger for split-operator MUX_2359_inst flow-through 
    process(IMA4_2360) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_2359_inst:flowthrough inputs: " & " BITSEL_u8_u1_2354_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_2354_wire) & " type_cast_2356_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2356_wire_constant) & " type_cast_2358_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2358_wire_constant) & " outputs:" & " IMA4_2360= "  & Convert_SLV_To_Hex_String(IMA4_2360));
      --
    end process; 
    -- flow-through select operator MUX_2359_inst
    IMA4_2360 <= type_cast_2356_wire_constant when (BITSEL_u8_u1_2354_wire(0) /=  '0') else type_cast_2358_wire_constant;
    -- logger for split-operator MUX_2369_inst flow-through 
    process(IMA5_2370) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_2369_inst:flowthrough inputs: " & " BITSEL_u8_u1_2364_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_2364_wire) & " type_cast_2366_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2366_wire_constant) & " type_cast_2368_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2368_wire_constant) & " outputs:" & " IMA5_2370= "  & Convert_SLV_To_Hex_String(IMA5_2370));
      --
    end process; 
    -- flow-through select operator MUX_2369_inst
    IMA5_2370 <= type_cast_2366_wire_constant when (BITSEL_u8_u1_2364_wire(0) /=  '0') else type_cast_2368_wire_constant;
    -- logger for split-operator MUX_2379_inst flow-through 
    process(IMA6_2380) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_2379_inst:flowthrough inputs: " & " BITSEL_u8_u1_2374_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_2374_wire) & " type_cast_2376_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2376_wire_constant) & " type_cast_2378_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2378_wire_constant) & " outputs:" & " IMA6_2380= "  & Convert_SLV_To_Hex_String(IMA6_2380));
      --
    end process; 
    -- flow-through select operator MUX_2379_inst
    IMA6_2380 <= type_cast_2376_wire_constant when (BITSEL_u8_u1_2374_wire(0) /=  '0') else type_cast_2378_wire_constant;
    -- logger for split-operator MUX_2389_inst flow-through 
    process(IMA7_2390) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_2389_inst:flowthrough inputs: " & " BITSEL_u8_u1_2384_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_2384_wire) & " type_cast_2386_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2386_wire_constant) & " type_cast_2388_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2388_wire_constant) & " outputs:" & " IMA7_2390= "  & Convert_SLV_To_Hex_String(IMA7_2390));
      --
    end process; 
    -- flow-through select operator MUX_2389_inst
    IMA7_2390 <= type_cast_2386_wire_constant when (BITSEL_u8_u1_2384_wire(0) /=  '0') else type_cast_2388_wire_constant;
    -- logger for split-operator MUX_2399_inst flow-through 
    process(IMA8_2400) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_2399_inst:flowthrough inputs: " & " BITSEL_u8_u1_2394_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_2394_wire) & " type_cast_2396_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2396_wire_constant) & " type_cast_2398_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2398_wire_constant) & " outputs:" & " IMA8_2400= "  & Convert_SLV_To_Hex_String(IMA8_2400));
      --
    end process; 
    -- flow-through select operator MUX_2399_inst
    IMA8_2400 <= type_cast_2396_wire_constant when (BITSEL_u8_u1_2394_wire(0) /=  '0') else type_cast_2398_wire_constant;
    -- logger for split-operator MUX_2409_inst flow-through 
    process(IMA9_2410) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_2409_inst:flowthrough inputs: " & " BITSEL_u8_u1_2404_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_2404_wire) & " type_cast_2406_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2406_wire_constant) & " type_cast_2408_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2408_wire_constant) & " outputs:" & " IMA9_2410= "  & Convert_SLV_To_Hex_String(IMA9_2410));
      --
    end process; 
    -- flow-through select operator MUX_2409_inst
    IMA9_2410 <= type_cast_2406_wire_constant when (BITSEL_u8_u1_2404_wire(0) /=  '0') else type_cast_2408_wire_constant;
    -- logger for split-operator MUX_2419_inst flow-through 
    process(IMA10_2420) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_2419_inst:flowthrough inputs: " & " BITSEL_u8_u1_2414_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_2414_wire) & " type_cast_2416_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2416_wire_constant) & " type_cast_2418_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2418_wire_constant) & " outputs:" & " IMA10_2420= "  & Convert_SLV_To_Hex_String(IMA10_2420));
      --
    end process; 
    -- flow-through select operator MUX_2419_inst
    IMA10_2420 <= type_cast_2416_wire_constant when (BITSEL_u8_u1_2414_wire(0) /=  '0') else type_cast_2418_wire_constant;
    -- logger for split-operator MUX_2429_inst flow-through 
    process(IMA11_2430) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_2429_inst:flowthrough inputs: " & " BITSEL_u8_u1_2424_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_2424_wire) & " type_cast_2426_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2426_wire_constant) & " type_cast_2428_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2428_wire_constant) & " outputs:" & " IMA11_2430= "  & Convert_SLV_To_Hex_String(IMA11_2430));
      --
    end process; 
    -- flow-through select operator MUX_2429_inst
    IMA11_2430 <= type_cast_2426_wire_constant when (BITSEL_u8_u1_2424_wire(0) /=  '0') else type_cast_2428_wire_constant;
    -- logger for split-operator MUX_2439_inst flow-through 
    process(IMA12_2440) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_2439_inst:flowthrough inputs: " & " BITSEL_u8_u1_2434_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_2434_wire) & " type_cast_2436_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2436_wire_constant) & " type_cast_2438_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2438_wire_constant) & " outputs:" & " IMA12_2440= "  & Convert_SLV_To_Hex_String(IMA12_2440));
      --
    end process; 
    -- flow-through select operator MUX_2439_inst
    IMA12_2440 <= type_cast_2436_wire_constant when (BITSEL_u8_u1_2434_wire(0) /=  '0') else type_cast_2438_wire_constant;
    -- logger for split-operator MUX_2449_inst flow-through 
    process(IMA13_2450) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_2449_inst:flowthrough inputs: " & " BITSEL_u8_u1_2444_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_2444_wire) & " type_cast_2446_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2446_wire_constant) & " type_cast_2448_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2448_wire_constant) & " outputs:" & " IMA13_2450= "  & Convert_SLV_To_Hex_String(IMA13_2450));
      --
    end process; 
    -- flow-through select operator MUX_2449_inst
    IMA13_2450 <= type_cast_2446_wire_constant when (BITSEL_u8_u1_2444_wire(0) /=  '0') else type_cast_2448_wire_constant;
    -- logger for split-operator MUX_2459_inst flow-through 
    process(IMA14_2460) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_2459_inst:flowthrough inputs: " & " BITSEL_u8_u1_2454_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_2454_wire) & " type_cast_2456_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2456_wire_constant) & " type_cast_2458_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2458_wire_constant) & " outputs:" & " IMA14_2460= "  & Convert_SLV_To_Hex_String(IMA14_2460));
      --
    end process; 
    -- flow-through select operator MUX_2459_inst
    IMA14_2460 <= type_cast_2456_wire_constant when (BITSEL_u8_u1_2454_wire(0) /=  '0') else type_cast_2458_wire_constant;
    -- logger for split-operator MUX_2469_inst flow-through 
    process(IMA15_2470) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_2469_inst:flowthrough inputs: " & " BITSEL_u8_u1_2464_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_2464_wire) & " type_cast_2466_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2466_wire_constant) & " type_cast_2468_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2468_wire_constant) & " outputs:" & " IMA15_2470= "  & Convert_SLV_To_Hex_String(IMA15_2470));
      --
    end process; 
    -- flow-through select operator MUX_2469_inst
    IMA15_2470 <= type_cast_2466_wire_constant when (BITSEL_u8_u1_2464_wire(0) /=  '0') else type_cast_2468_wire_constant;
    -- logger for split-operator MUX_2479_inst flow-through 
    process(IMA16_2480) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_2479_inst:flowthrough inputs: " & " BITSEL_u8_u1_2474_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_2474_wire) & " type_cast_2476_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2476_wire_constant) & " type_cast_2478_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2478_wire_constant) & " outputs:" & " IMA16_2480= "  & Convert_SLV_To_Hex_String(IMA16_2480));
      --
    end process; 
    -- flow-through select operator MUX_2479_inst
    IMA16_2480 <= type_cast_2476_wire_constant when (BITSEL_u8_u1_2474_wire(0) /=  '0') else type_cast_2478_wire_constant;
    -- logger for split-operator MUX_2489_inst flow-through 
    process(IMA17_2490) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_2489_inst:flowthrough inputs: " & " BITSEL_u8_u1_2484_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_2484_wire) & " type_cast_2486_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2486_wire_constant) & " type_cast_2488_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2488_wire_constant) & " outputs:" & " IMA17_2490= "  & Convert_SLV_To_Hex_String(IMA17_2490));
      --
    end process; 
    -- flow-through select operator MUX_2489_inst
    IMA17_2490 <= type_cast_2486_wire_constant when (BITSEL_u8_u1_2484_wire(0) /=  '0') else type_cast_2488_wire_constant;
    -- logger for split-operator MUX_2499_inst flow-through 
    process(IMA18_2500) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_2499_inst:flowthrough inputs: " & " BITSEL_u8_u1_2494_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_2494_wire) & " type_cast_2496_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2496_wire_constant) & " type_cast_2498_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2498_wire_constant) & " outputs:" & " IMA18_2500= "  & Convert_SLV_To_Hex_String(IMA18_2500));
      --
    end process; 
    -- flow-through select operator MUX_2499_inst
    IMA18_2500 <= type_cast_2496_wire_constant when (BITSEL_u8_u1_2494_wire(0) /=  '0') else type_cast_2498_wire_constant;
    -- logger for split-operator MUX_2509_inst flow-through 
    process(IMA19_2510) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_2509_inst:flowthrough inputs: " & " BITSEL_u8_u1_2504_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_2504_wire) & " type_cast_2506_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2506_wire_constant) & " type_cast_2508_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2508_wire_constant) & " outputs:" & " IMA19_2510= "  & Convert_SLV_To_Hex_String(IMA19_2510));
      --
    end process; 
    -- flow-through select operator MUX_2509_inst
    IMA19_2510 <= type_cast_2506_wire_constant when (BITSEL_u8_u1_2504_wire(0) /=  '0') else type_cast_2508_wire_constant;
    -- logger for split-operator MUX_2519_inst flow-through 
    process(IMA20_2520) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_2519_inst:flowthrough inputs: " & " BITSEL_u8_u1_2514_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_2514_wire) & " type_cast_2516_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2516_wire_constant) & " type_cast_2518_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2518_wire_constant) & " outputs:" & " IMA20_2520= "  & Convert_SLV_To_Hex_String(IMA20_2520));
      --
    end process; 
    -- flow-through select operator MUX_2519_inst
    IMA20_2520 <= type_cast_2516_wire_constant when (BITSEL_u8_u1_2514_wire(0) /=  '0') else type_cast_2518_wire_constant;
    -- logger for split-operator MUX_2529_inst flow-through 
    process(IMA21_2530) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_2529_inst:flowthrough inputs: " & " BITSEL_u8_u1_2524_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_2524_wire) & " type_cast_2526_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2526_wire_constant) & " type_cast_2528_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2528_wire_constant) & " outputs:" & " IMA21_2530= "  & Convert_SLV_To_Hex_String(IMA21_2530));
      --
    end process; 
    -- flow-through select operator MUX_2529_inst
    IMA21_2530 <= type_cast_2526_wire_constant when (BITSEL_u8_u1_2524_wire(0) /=  '0') else type_cast_2528_wire_constant;
    -- logger for split-operator MUX_2539_inst flow-through 
    process(IMA22_2540) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_2539_inst:flowthrough inputs: " & " BITSEL_u8_u1_2534_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_2534_wire) & " type_cast_2536_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2536_wire_constant) & " type_cast_2538_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2538_wire_constant) & " outputs:" & " IMA22_2540= "  & Convert_SLV_To_Hex_String(IMA22_2540));
      --
    end process; 
    -- flow-through select operator MUX_2539_inst
    IMA22_2540 <= type_cast_2536_wire_constant when (BITSEL_u8_u1_2534_wire(0) /=  '0') else type_cast_2538_wire_constant;
    -- logger for split-operator MUX_2549_inst flow-through 
    process(IMA23_2550) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_2549_inst:flowthrough inputs: " & " BITSEL_u8_u1_2544_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_2544_wire) & " type_cast_2546_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2546_wire_constant) & " type_cast_2548_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2548_wire_constant) & " outputs:" & " IMA23_2550= "  & Convert_SLV_To_Hex_String(IMA23_2550));
      --
    end process; 
    -- flow-through select operator MUX_2549_inst
    IMA23_2550 <= type_cast_2546_wire_constant when (BITSEL_u8_u1_2544_wire(0) /=  '0') else type_cast_2548_wire_constant;
    -- logger for split-operator MUX_2559_inst flow-through 
    process(IMA24_2560) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_2559_inst:flowthrough inputs: " & " BITSEL_u8_u1_2554_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_2554_wire) & " type_cast_2556_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2556_wire_constant) & " type_cast_2558_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2558_wire_constant) & " outputs:" & " IMA24_2560= "  & Convert_SLV_To_Hex_String(IMA24_2560));
      --
    end process; 
    -- flow-through select operator MUX_2559_inst
    IMA24_2560 <= type_cast_2556_wire_constant when (BITSEL_u8_u1_2554_wire(0) /=  '0') else type_cast_2558_wire_constant;
    -- logger for split-operator MUX_2569_inst flow-through 
    process(IMA25_2570) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_2569_inst:flowthrough inputs: " & " BITSEL_u8_u1_2564_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_2564_wire) & " type_cast_2566_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2566_wire_constant) & " type_cast_2568_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2568_wire_constant) & " outputs:" & " IMA25_2570= "  & Convert_SLV_To_Hex_String(IMA25_2570));
      --
    end process; 
    -- flow-through select operator MUX_2569_inst
    IMA25_2570 <= type_cast_2566_wire_constant when (BITSEL_u8_u1_2564_wire(0) /=  '0') else type_cast_2568_wire_constant;
    -- logger for split-operator MUX_2579_inst flow-through 
    process(IMA26_2580) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_2579_inst:flowthrough inputs: " & " BITSEL_u8_u1_2574_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_2574_wire) & " type_cast_2576_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2576_wire_constant) & " type_cast_2578_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2578_wire_constant) & " outputs:" & " IMA26_2580= "  & Convert_SLV_To_Hex_String(IMA26_2580));
      --
    end process; 
    -- flow-through select operator MUX_2579_inst
    IMA26_2580 <= type_cast_2576_wire_constant when (BITSEL_u8_u1_2574_wire(0) /=  '0') else type_cast_2578_wire_constant;
    -- logger for split-operator MUX_2589_inst flow-through 
    process(IMA27_2590) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_2589_inst:flowthrough inputs: " & " BITSEL_u8_u1_2584_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_2584_wire) & " type_cast_2586_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2586_wire_constant) & " type_cast_2588_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2588_wire_constant) & " outputs:" & " IMA27_2590= "  & Convert_SLV_To_Hex_String(IMA27_2590));
      --
    end process; 
    -- flow-through select operator MUX_2589_inst
    IMA27_2590 <= type_cast_2586_wire_constant when (BITSEL_u8_u1_2584_wire(0) /=  '0') else type_cast_2588_wire_constant;
    -- logger for split-operator MUX_2599_inst flow-through 
    process(IMA28_2600) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_2599_inst:flowthrough inputs: " & " BITSEL_u8_u1_2594_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_2594_wire) & " type_cast_2596_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2596_wire_constant) & " type_cast_2598_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2598_wire_constant) & " outputs:" & " IMA28_2600= "  & Convert_SLV_To_Hex_String(IMA28_2600));
      --
    end process; 
    -- flow-through select operator MUX_2599_inst
    IMA28_2600 <= type_cast_2596_wire_constant when (BITSEL_u8_u1_2594_wire(0) /=  '0') else type_cast_2598_wire_constant;
    -- logger for split-operator MUX_2609_inst flow-through 
    process(IMA29_2610) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_2609_inst:flowthrough inputs: " & " BITSEL_u8_u1_2604_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_2604_wire) & " type_cast_2606_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2606_wire_constant) & " type_cast_2608_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2608_wire_constant) & " outputs:" & " IMA29_2610= "  & Convert_SLV_To_Hex_String(IMA29_2610));
      --
    end process; 
    -- flow-through select operator MUX_2609_inst
    IMA29_2610 <= type_cast_2606_wire_constant when (BITSEL_u8_u1_2604_wire(0) /=  '0') else type_cast_2608_wire_constant;
    -- logger for split-operator MUX_2619_inst flow-through 
    process(IMA30_2620) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_2619_inst:flowthrough inputs: " & " BITSEL_u8_u1_2614_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_2614_wire) & " type_cast_2616_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2616_wire_constant) & " type_cast_2618_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2618_wire_constant) & " outputs:" & " IMA30_2620= "  & Convert_SLV_To_Hex_String(IMA30_2620));
      --
    end process; 
    -- flow-through select operator MUX_2619_inst
    IMA30_2620 <= type_cast_2616_wire_constant when (BITSEL_u8_u1_2614_wire(0) /=  '0') else type_cast_2618_wire_constant;
    -- logger for split-operator MUX_2629_inst flow-through 
    process(IMA31_2630) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_2629_inst:flowthrough inputs: " & " BITSEL_u8_u1_2624_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_2624_wire) & " type_cast_2626_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2626_wire_constant) & " type_cast_2628_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2628_wire_constant) & " outputs:" & " IMA31_2630= "  & Convert_SLV_To_Hex_String(IMA31_2630));
      --
    end process; 
    -- flow-through select operator MUX_2629_inst
    IMA31_2630 <= type_cast_2626_wire_constant when (BITSEL_u8_u1_2624_wire(0) /=  '0') else type_cast_2628_wire_constant;
    -- logger for split-operator MUX_2639_inst flow-through 
    process(IMA32_2640) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_2639_inst:flowthrough inputs: " & " BITSEL_u8_u1_2634_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_2634_wire) & " type_cast_2636_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2636_wire_constant) & " type_cast_2638_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2638_wire_constant) & " outputs:" & " IMA32_2640= "  & Convert_SLV_To_Hex_String(IMA32_2640));
      --
    end process; 
    -- flow-through select operator MUX_2639_inst
    IMA32_2640 <= type_cast_2636_wire_constant when (BITSEL_u8_u1_2634_wire(0) /=  '0') else type_cast_2638_wire_constant;
    -- logger for split-operator MUX_2649_inst flow-through 
    process(IMA33_2650) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_2649_inst:flowthrough inputs: " & " BITSEL_u8_u1_2644_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_2644_wire) & " type_cast_2646_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2646_wire_constant) & " type_cast_2648_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2648_wire_constant) & " outputs:" & " IMA33_2650= "  & Convert_SLV_To_Hex_String(IMA33_2650));
      --
    end process; 
    -- flow-through select operator MUX_2649_inst
    IMA33_2650 <= type_cast_2646_wire_constant when (BITSEL_u8_u1_2644_wire(0) /=  '0') else type_cast_2648_wire_constant;
    -- logger for split-operator MUX_2659_inst flow-through 
    process(IMA34_2660) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_2659_inst:flowthrough inputs: " & " BITSEL_u8_u1_2654_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_2654_wire) & " type_cast_2656_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2656_wire_constant) & " type_cast_2658_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2658_wire_constant) & " outputs:" & " IMA34_2660= "  & Convert_SLV_To_Hex_String(IMA34_2660));
      --
    end process; 
    -- flow-through select operator MUX_2659_inst
    IMA34_2660 <= type_cast_2656_wire_constant when (BITSEL_u8_u1_2654_wire(0) /=  '0') else type_cast_2658_wire_constant;
    -- logger for split-operator MUX_2669_inst flow-through 
    process(IMA35_2670) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_2669_inst:flowthrough inputs: " & " BITSEL_u8_u1_2664_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_2664_wire) & " type_cast_2666_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2666_wire_constant) & " type_cast_2668_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2668_wire_constant) & " outputs:" & " IMA35_2670= "  & Convert_SLV_To_Hex_String(IMA35_2670));
      --
    end process; 
    -- flow-through select operator MUX_2669_inst
    IMA35_2670 <= type_cast_2666_wire_constant when (BITSEL_u8_u1_2664_wire(0) /=  '0') else type_cast_2668_wire_constant;
    -- logger for split-operator MUX_2679_inst flow-through 
    process(IMA36_2680) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_2679_inst:flowthrough inputs: " & " BITSEL_u8_u1_2674_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_2674_wire) & " type_cast_2676_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2676_wire_constant) & " type_cast_2678_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2678_wire_constant) & " outputs:" & " IMA36_2680= "  & Convert_SLV_To_Hex_String(IMA36_2680));
      --
    end process; 
    -- flow-through select operator MUX_2679_inst
    IMA36_2680 <= type_cast_2676_wire_constant when (BITSEL_u8_u1_2674_wire(0) /=  '0') else type_cast_2678_wire_constant;
    -- logger for split-operator MUX_2689_inst flow-through 
    process(IMA37_2690) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_2689_inst:flowthrough inputs: " & " BITSEL_u8_u1_2684_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_2684_wire) & " type_cast_2686_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2686_wire_constant) & " type_cast_2688_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2688_wire_constant) & " outputs:" & " IMA37_2690= "  & Convert_SLV_To_Hex_String(IMA37_2690));
      --
    end process; 
    -- flow-through select operator MUX_2689_inst
    IMA37_2690 <= type_cast_2686_wire_constant when (BITSEL_u8_u1_2684_wire(0) /=  '0') else type_cast_2688_wire_constant;
    -- logger for split-operator MUX_2699_inst flow-through 
    process(IMA38_2700) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_2699_inst:flowthrough inputs: " & " BITSEL_u8_u1_2694_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_2694_wire) & " type_cast_2696_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2696_wire_constant) & " type_cast_2698_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2698_wire_constant) & " outputs:" & " IMA38_2700= "  & Convert_SLV_To_Hex_String(IMA38_2700));
      --
    end process; 
    -- flow-through select operator MUX_2699_inst
    IMA38_2700 <= type_cast_2696_wire_constant when (BITSEL_u8_u1_2694_wire(0) /=  '0') else type_cast_2698_wire_constant;
    -- logger for split-operator MUX_2709_inst flow-through 
    process(IMA39_2710) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_2709_inst:flowthrough inputs: " & " BITSEL_u8_u1_2704_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_2704_wire) & " type_cast_2706_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2706_wire_constant) & " type_cast_2708_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2708_wire_constant) & " outputs:" & " IMA39_2710= "  & Convert_SLV_To_Hex_String(IMA39_2710));
      --
    end process; 
    -- flow-through select operator MUX_2709_inst
    IMA39_2710 <= type_cast_2706_wire_constant when (BITSEL_u8_u1_2704_wire(0) /=  '0') else type_cast_2708_wire_constant;
    -- logger for split-operator MUX_2719_inst flow-through 
    process(IMA40_2720) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_2719_inst:flowthrough inputs: " & " BITSEL_u8_u1_2714_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_2714_wire) & " type_cast_2716_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2716_wire_constant) & " type_cast_2718_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2718_wire_constant) & " outputs:" & " IMA40_2720= "  & Convert_SLV_To_Hex_String(IMA40_2720));
      --
    end process; 
    -- flow-through select operator MUX_2719_inst
    IMA40_2720 <= type_cast_2716_wire_constant when (BITSEL_u8_u1_2714_wire(0) /=  '0') else type_cast_2718_wire_constant;
    -- logger for split-operator MUX_2729_inst flow-through 
    process(IMA41_2730) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_2729_inst:flowthrough inputs: " & " BITSEL_u8_u1_2724_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_2724_wire) & " type_cast_2726_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2726_wire_constant) & " type_cast_2728_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2728_wire_constant) & " outputs:" & " IMA41_2730= "  & Convert_SLV_To_Hex_String(IMA41_2730));
      --
    end process; 
    -- flow-through select operator MUX_2729_inst
    IMA41_2730 <= type_cast_2726_wire_constant when (BITSEL_u8_u1_2724_wire(0) /=  '0') else type_cast_2728_wire_constant;
    -- logger for split-operator MUX_2739_inst flow-through 
    process(IMA42_2740) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_2739_inst:flowthrough inputs: " & " BITSEL_u8_u1_2734_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_2734_wire) & " type_cast_2736_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2736_wire_constant) & " type_cast_2738_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2738_wire_constant) & " outputs:" & " IMA42_2740= "  & Convert_SLV_To_Hex_String(IMA42_2740));
      --
    end process; 
    -- flow-through select operator MUX_2739_inst
    IMA42_2740 <= type_cast_2736_wire_constant when (BITSEL_u8_u1_2734_wire(0) /=  '0') else type_cast_2738_wire_constant;
    -- logger for split-operator MUX_2749_inst flow-through 
    process(IMA43_2750) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_2749_inst:flowthrough inputs: " & " BITSEL_u8_u1_2744_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_2744_wire) & " type_cast_2746_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2746_wire_constant) & " type_cast_2748_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2748_wire_constant) & " outputs:" & " IMA43_2750= "  & Convert_SLV_To_Hex_String(IMA43_2750));
      --
    end process; 
    -- flow-through select operator MUX_2749_inst
    IMA43_2750 <= type_cast_2746_wire_constant when (BITSEL_u8_u1_2744_wire(0) /=  '0') else type_cast_2748_wire_constant;
    -- logger for split-operator MUX_2759_inst flow-through 
    process(IMA44_2760) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_2759_inst:flowthrough inputs: " & " BITSEL_u8_u1_2754_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_2754_wire) & " type_cast_2756_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2756_wire_constant) & " type_cast_2758_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2758_wire_constant) & " outputs:" & " IMA44_2760= "  & Convert_SLV_To_Hex_String(IMA44_2760));
      --
    end process; 
    -- flow-through select operator MUX_2759_inst
    IMA44_2760 <= type_cast_2756_wire_constant when (BITSEL_u8_u1_2754_wire(0) /=  '0') else type_cast_2758_wire_constant;
    -- logger for split-operator MUX_2769_inst flow-through 
    process(IMA45_2770) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_2769_inst:flowthrough inputs: " & " BITSEL_u8_u1_2764_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_2764_wire) & " type_cast_2766_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2766_wire_constant) & " type_cast_2768_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2768_wire_constant) & " outputs:" & " IMA45_2770= "  & Convert_SLV_To_Hex_String(IMA45_2770));
      --
    end process; 
    -- flow-through select operator MUX_2769_inst
    IMA45_2770 <= type_cast_2766_wire_constant when (BITSEL_u8_u1_2764_wire(0) /=  '0') else type_cast_2768_wire_constant;
    -- logger for split-operator MUX_2779_inst flow-through 
    process(IMA46_2780) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_2779_inst:flowthrough inputs: " & " BITSEL_u8_u1_2774_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_2774_wire) & " type_cast_2776_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2776_wire_constant) & " type_cast_2778_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2778_wire_constant) & " outputs:" & " IMA46_2780= "  & Convert_SLV_To_Hex_String(IMA46_2780));
      --
    end process; 
    -- flow-through select operator MUX_2779_inst
    IMA46_2780 <= type_cast_2776_wire_constant when (BITSEL_u8_u1_2774_wire(0) /=  '0') else type_cast_2778_wire_constant;
    -- logger for split-operator MUX_2789_inst flow-through 
    process(IMA47_2790) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_2789_inst:flowthrough inputs: " & " BITSEL_u8_u1_2784_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_2784_wire) & " type_cast_2786_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2786_wire_constant) & " type_cast_2788_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2788_wire_constant) & " outputs:" & " IMA47_2790= "  & Convert_SLV_To_Hex_String(IMA47_2790));
      --
    end process; 
    -- flow-through select operator MUX_2789_inst
    IMA47_2790 <= type_cast_2786_wire_constant when (BITSEL_u8_u1_2784_wire(0) /=  '0') else type_cast_2788_wire_constant;
    -- logger for split-operator MUX_2799_inst flow-through 
    process(IMA48_2800) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_2799_inst:flowthrough inputs: " & " BITSEL_u8_u1_2794_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_2794_wire) & " type_cast_2796_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2796_wire_constant) & " type_cast_2798_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2798_wire_constant) & " outputs:" & " IMA48_2800= "  & Convert_SLV_To_Hex_String(IMA48_2800));
      --
    end process; 
    -- flow-through select operator MUX_2799_inst
    IMA48_2800 <= type_cast_2796_wire_constant when (BITSEL_u8_u1_2794_wire(0) /=  '0') else type_cast_2798_wire_constant;
    -- logger for split-operator MUX_2809_inst flow-through 
    process(IMA49_2810) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_2809_inst:flowthrough inputs: " & " BITSEL_u8_u1_2804_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_2804_wire) & " type_cast_2806_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2806_wire_constant) & " type_cast_2808_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2808_wire_constant) & " outputs:" & " IMA49_2810= "  & Convert_SLV_To_Hex_String(IMA49_2810));
      --
    end process; 
    -- flow-through select operator MUX_2809_inst
    IMA49_2810 <= type_cast_2806_wire_constant when (BITSEL_u8_u1_2804_wire(0) /=  '0') else type_cast_2808_wire_constant;
    -- logger for split-operator MUX_2819_inst flow-through 
    process(IMA50_2820) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_2819_inst:flowthrough inputs: " & " BITSEL_u8_u1_2814_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_2814_wire) & " type_cast_2816_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2816_wire_constant) & " type_cast_2818_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2818_wire_constant) & " outputs:" & " IMA50_2820= "  & Convert_SLV_To_Hex_String(IMA50_2820));
      --
    end process; 
    -- flow-through select operator MUX_2819_inst
    IMA50_2820 <= type_cast_2816_wire_constant when (BITSEL_u8_u1_2814_wire(0) /=  '0') else type_cast_2818_wire_constant;
    -- logger for split-operator MUX_2829_inst flow-through 
    process(IMA51_2830) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_2829_inst:flowthrough inputs: " & " BITSEL_u8_u1_2824_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_2824_wire) & " type_cast_2826_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2826_wire_constant) & " type_cast_2828_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2828_wire_constant) & " outputs:" & " IMA51_2830= "  & Convert_SLV_To_Hex_String(IMA51_2830));
      --
    end process; 
    -- flow-through select operator MUX_2829_inst
    IMA51_2830 <= type_cast_2826_wire_constant when (BITSEL_u8_u1_2824_wire(0) /=  '0') else type_cast_2828_wire_constant;
    -- logger for split-operator MUX_2839_inst flow-through 
    process(IMA52_2840) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_2839_inst:flowthrough inputs: " & " BITSEL_u8_u1_2834_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_2834_wire) & " type_cast_2836_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2836_wire_constant) & " type_cast_2838_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2838_wire_constant) & " outputs:" & " IMA52_2840= "  & Convert_SLV_To_Hex_String(IMA52_2840));
      --
    end process; 
    -- flow-through select operator MUX_2839_inst
    IMA52_2840 <= type_cast_2836_wire_constant when (BITSEL_u8_u1_2834_wire(0) /=  '0') else type_cast_2838_wire_constant;
    -- logger for split-operator MUX_2849_inst flow-through 
    process(IMA53_2850) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_2849_inst:flowthrough inputs: " & " BITSEL_u8_u1_2844_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_2844_wire) & " type_cast_2846_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2846_wire_constant) & " type_cast_2848_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2848_wire_constant) & " outputs:" & " IMA53_2850= "  & Convert_SLV_To_Hex_String(IMA53_2850));
      --
    end process; 
    -- flow-through select operator MUX_2849_inst
    IMA53_2850 <= type_cast_2846_wire_constant when (BITSEL_u8_u1_2844_wire(0) /=  '0') else type_cast_2848_wire_constant;
    -- logger for split-operator MUX_2859_inst flow-through 
    process(IMA54_2860) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_2859_inst:flowthrough inputs: " & " BITSEL_u8_u1_2854_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_2854_wire) & " type_cast_2856_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2856_wire_constant) & " type_cast_2858_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2858_wire_constant) & " outputs:" & " IMA54_2860= "  & Convert_SLV_To_Hex_String(IMA54_2860));
      --
    end process; 
    -- flow-through select operator MUX_2859_inst
    IMA54_2860 <= type_cast_2856_wire_constant when (BITSEL_u8_u1_2854_wire(0) /=  '0') else type_cast_2858_wire_constant;
    -- logger for split-operator MUX_2869_inst flow-through 
    process(IMA55_2870) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_2869_inst:flowthrough inputs: " & " BITSEL_u8_u1_2864_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_2864_wire) & " type_cast_2866_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2866_wire_constant) & " type_cast_2868_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2868_wire_constant) & " outputs:" & " IMA55_2870= "  & Convert_SLV_To_Hex_String(IMA55_2870));
      --
    end process; 
    -- flow-through select operator MUX_2869_inst
    IMA55_2870 <= type_cast_2866_wire_constant when (BITSEL_u8_u1_2864_wire(0) /=  '0') else type_cast_2868_wire_constant;
    -- logger for split-operator MUX_2879_inst flow-through 
    process(IMA56_2880) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_2879_inst:flowthrough inputs: " & " BITSEL_u8_u1_2874_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_2874_wire) & " type_cast_2876_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2876_wire_constant) & " type_cast_2878_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2878_wire_constant) & " outputs:" & " IMA56_2880= "  & Convert_SLV_To_Hex_String(IMA56_2880));
      --
    end process; 
    -- flow-through select operator MUX_2879_inst
    IMA56_2880 <= type_cast_2876_wire_constant when (BITSEL_u8_u1_2874_wire(0) /=  '0') else type_cast_2878_wire_constant;
    -- logger for split-operator MUX_2889_inst flow-through 
    process(IMA57_2890) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_2889_inst:flowthrough inputs: " & " BITSEL_u8_u1_2884_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_2884_wire) & " type_cast_2886_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2886_wire_constant) & " type_cast_2888_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2888_wire_constant) & " outputs:" & " IMA57_2890= "  & Convert_SLV_To_Hex_String(IMA57_2890));
      --
    end process; 
    -- flow-through select operator MUX_2889_inst
    IMA57_2890 <= type_cast_2886_wire_constant when (BITSEL_u8_u1_2884_wire(0) /=  '0') else type_cast_2888_wire_constant;
    -- logger for split-operator MUX_2899_inst flow-through 
    process(IMA58_2900) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_2899_inst:flowthrough inputs: " & " BITSEL_u8_u1_2894_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_2894_wire) & " type_cast_2896_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2896_wire_constant) & " type_cast_2898_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2898_wire_constant) & " outputs:" & " IMA58_2900= "  & Convert_SLV_To_Hex_String(IMA58_2900));
      --
    end process; 
    -- flow-through select operator MUX_2899_inst
    IMA58_2900 <= type_cast_2896_wire_constant when (BITSEL_u8_u1_2894_wire(0) /=  '0') else type_cast_2898_wire_constant;
    -- logger for split-operator MUX_2909_inst flow-through 
    process(IMA59_2910) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_2909_inst:flowthrough inputs: " & " BITSEL_u8_u1_2904_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_2904_wire) & " type_cast_2906_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2906_wire_constant) & " type_cast_2908_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2908_wire_constant) & " outputs:" & " IMA59_2910= "  & Convert_SLV_To_Hex_String(IMA59_2910));
      --
    end process; 
    -- flow-through select operator MUX_2909_inst
    IMA59_2910 <= type_cast_2906_wire_constant when (BITSEL_u8_u1_2904_wire(0) /=  '0') else type_cast_2908_wire_constant;
    -- logger for split-operator MUX_2919_inst flow-through 
    process(IMA60_2920) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_2919_inst:flowthrough inputs: " & " BITSEL_u8_u1_2914_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_2914_wire) & " type_cast_2916_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2916_wire_constant) & " type_cast_2918_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2918_wire_constant) & " outputs:" & " IMA60_2920= "  & Convert_SLV_To_Hex_String(IMA60_2920));
      --
    end process; 
    -- flow-through select operator MUX_2919_inst
    IMA60_2920 <= type_cast_2916_wire_constant when (BITSEL_u8_u1_2914_wire(0) /=  '0') else type_cast_2918_wire_constant;
    -- logger for split-operator MUX_2929_inst flow-through 
    process(IMA61_2930) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_2929_inst:flowthrough inputs: " & " BITSEL_u8_u1_2924_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_2924_wire) & " type_cast_2926_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2926_wire_constant) & " type_cast_2928_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2928_wire_constant) & " outputs:" & " IMA61_2930= "  & Convert_SLV_To_Hex_String(IMA61_2930));
      --
    end process; 
    -- flow-through select operator MUX_2929_inst
    IMA61_2930 <= type_cast_2926_wire_constant when (BITSEL_u8_u1_2924_wire(0) /=  '0') else type_cast_2928_wire_constant;
    -- logger for split-operator MUX_2939_inst flow-through 
    process(IMA62_2940) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_2939_inst:flowthrough inputs: " & " BITSEL_u8_u1_2934_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_2934_wire) & " type_cast_2936_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2936_wire_constant) & " type_cast_2938_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2938_wire_constant) & " outputs:" & " IMA62_2940= "  & Convert_SLV_To_Hex_String(IMA62_2940));
      --
    end process; 
    -- flow-through select operator MUX_2939_inst
    IMA62_2940 <= type_cast_2936_wire_constant when (BITSEL_u8_u1_2934_wire(0) /=  '0') else type_cast_2938_wire_constant;
    -- logger for split-operator MUX_2949_inst flow-through 
    process(IMA63_2950) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_2949_inst:flowthrough inputs: " & " BITSEL_u8_u1_2944_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_2944_wire) & " type_cast_2946_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2946_wire_constant) & " type_cast_2948_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2948_wire_constant) & " outputs:" & " IMA63_2950= "  & Convert_SLV_To_Hex_String(IMA63_2950));
      --
    end process; 
    -- flow-through select operator MUX_2949_inst
    IMA63_2950 <= type_cast_2946_wire_constant when (BITSEL_u8_u1_2944_wire(0) /=  '0') else type_cast_2948_wire_constant;
    -- logger for split-operator MUX_2959_inst flow-through 
    process(IMA64_2960) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_2959_inst:flowthrough inputs: " & " BITSEL_u8_u1_2954_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_2954_wire) & " type_cast_2956_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2956_wire_constant) & " type_cast_2958_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2958_wire_constant) & " outputs:" & " IMA64_2960= "  & Convert_SLV_To_Hex_String(IMA64_2960));
      --
    end process; 
    -- flow-through select operator MUX_2959_inst
    IMA64_2960 <= type_cast_2956_wire_constant when (BITSEL_u8_u1_2954_wire(0) /=  '0') else type_cast_2958_wire_constant;
    -- logger for split-operator MUX_2969_inst flow-through 
    process(IMA65_2970) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_2969_inst:flowthrough inputs: " & " BITSEL_u8_u1_2964_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_2964_wire) & " type_cast_2966_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2966_wire_constant) & " type_cast_2968_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2968_wire_constant) & " outputs:" & " IMA65_2970= "  & Convert_SLV_To_Hex_String(IMA65_2970));
      --
    end process; 
    -- flow-through select operator MUX_2969_inst
    IMA65_2970 <= type_cast_2966_wire_constant when (BITSEL_u8_u1_2964_wire(0) /=  '0') else type_cast_2968_wire_constant;
    -- logger for split-operator MUX_2979_inst flow-through 
    process(IMA66_2980) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_2979_inst:flowthrough inputs: " & " BITSEL_u8_u1_2974_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_2974_wire) & " type_cast_2976_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2976_wire_constant) & " type_cast_2978_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2978_wire_constant) & " outputs:" & " IMA66_2980= "  & Convert_SLV_To_Hex_String(IMA66_2980));
      --
    end process; 
    -- flow-through select operator MUX_2979_inst
    IMA66_2980 <= type_cast_2976_wire_constant when (BITSEL_u8_u1_2974_wire(0) /=  '0') else type_cast_2978_wire_constant;
    -- logger for split-operator MUX_2989_inst flow-through 
    process(IMA67_2990) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_2989_inst:flowthrough inputs: " & " BITSEL_u8_u1_2984_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_2984_wire) & " type_cast_2986_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2986_wire_constant) & " type_cast_2988_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2988_wire_constant) & " outputs:" & " IMA67_2990= "  & Convert_SLV_To_Hex_String(IMA67_2990));
      --
    end process; 
    -- flow-through select operator MUX_2989_inst
    IMA67_2990 <= type_cast_2986_wire_constant when (BITSEL_u8_u1_2984_wire(0) /=  '0') else type_cast_2988_wire_constant;
    -- logger for split-operator MUX_2999_inst flow-through 
    process(IMA68_3000) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_2999_inst:flowthrough inputs: " & " BITSEL_u8_u1_2994_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_2994_wire) & " type_cast_2996_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2996_wire_constant) & " type_cast_2998_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2998_wire_constant) & " outputs:" & " IMA68_3000= "  & Convert_SLV_To_Hex_String(IMA68_3000));
      --
    end process; 
    -- flow-through select operator MUX_2999_inst
    IMA68_3000 <= type_cast_2996_wire_constant when (BITSEL_u8_u1_2994_wire(0) /=  '0') else type_cast_2998_wire_constant;
    -- logger for split-operator MUX_3009_inst flow-through 
    process(IMA69_3010) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3009_inst:flowthrough inputs: " & " BITSEL_u8_u1_3004_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3004_wire) & " type_cast_3006_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3006_wire_constant) & " type_cast_3008_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3008_wire_constant) & " outputs:" & " IMA69_3010= "  & Convert_SLV_To_Hex_String(IMA69_3010));
      --
    end process; 
    -- flow-through select operator MUX_3009_inst
    IMA69_3010 <= type_cast_3006_wire_constant when (BITSEL_u8_u1_3004_wire(0) /=  '0') else type_cast_3008_wire_constant;
    -- logger for split-operator MUX_3019_inst flow-through 
    process(IMA70_3020) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3019_inst:flowthrough inputs: " & " BITSEL_u8_u1_3014_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3014_wire) & " type_cast_3016_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3016_wire_constant) & " type_cast_3018_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3018_wire_constant) & " outputs:" & " IMA70_3020= "  & Convert_SLV_To_Hex_String(IMA70_3020));
      --
    end process; 
    -- flow-through select operator MUX_3019_inst
    IMA70_3020 <= type_cast_3016_wire_constant when (BITSEL_u8_u1_3014_wire(0) /=  '0') else type_cast_3018_wire_constant;
    -- logger for split-operator MUX_3029_inst flow-through 
    process(IMA71_3030) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3029_inst:flowthrough inputs: " & " BITSEL_u8_u1_3024_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3024_wire) & " type_cast_3026_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3026_wire_constant) & " type_cast_3028_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3028_wire_constant) & " outputs:" & " IMA71_3030= "  & Convert_SLV_To_Hex_String(IMA71_3030));
      --
    end process; 
    -- flow-through select operator MUX_3029_inst
    IMA71_3030 <= type_cast_3026_wire_constant when (BITSEL_u8_u1_3024_wire(0) /=  '0') else type_cast_3028_wire_constant;
    -- logger for split-operator MUX_3039_inst flow-through 
    process(IMA72_3040) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3039_inst:flowthrough inputs: " & " BITSEL_u8_u1_3034_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3034_wire) & " type_cast_3036_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3036_wire_constant) & " type_cast_3038_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3038_wire_constant) & " outputs:" & " IMA72_3040= "  & Convert_SLV_To_Hex_String(IMA72_3040));
      --
    end process; 
    -- flow-through select operator MUX_3039_inst
    IMA72_3040 <= type_cast_3036_wire_constant when (BITSEL_u8_u1_3034_wire(0) /=  '0') else type_cast_3038_wire_constant;
    -- logger for split-operator MUX_3049_inst flow-through 
    process(IMA73_3050) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3049_inst:flowthrough inputs: " & " BITSEL_u8_u1_3044_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3044_wire) & " type_cast_3046_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3046_wire_constant) & " type_cast_3048_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3048_wire_constant) & " outputs:" & " IMA73_3050= "  & Convert_SLV_To_Hex_String(IMA73_3050));
      --
    end process; 
    -- flow-through select operator MUX_3049_inst
    IMA73_3050 <= type_cast_3046_wire_constant when (BITSEL_u8_u1_3044_wire(0) /=  '0') else type_cast_3048_wire_constant;
    -- logger for split-operator MUX_3059_inst flow-through 
    process(IMA74_3060) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3059_inst:flowthrough inputs: " & " BITSEL_u8_u1_3054_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3054_wire) & " type_cast_3056_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3056_wire_constant) & " type_cast_3058_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3058_wire_constant) & " outputs:" & " IMA74_3060= "  & Convert_SLV_To_Hex_String(IMA74_3060));
      --
    end process; 
    -- flow-through select operator MUX_3059_inst
    IMA74_3060 <= type_cast_3056_wire_constant when (BITSEL_u8_u1_3054_wire(0) /=  '0') else type_cast_3058_wire_constant;
    -- logger for split-operator MUX_3069_inst flow-through 
    process(IMA75_3070) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3069_inst:flowthrough inputs: " & " BITSEL_u8_u1_3064_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3064_wire) & " type_cast_3066_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3066_wire_constant) & " type_cast_3068_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3068_wire_constant) & " outputs:" & " IMA75_3070= "  & Convert_SLV_To_Hex_String(IMA75_3070));
      --
    end process; 
    -- flow-through select operator MUX_3069_inst
    IMA75_3070 <= type_cast_3066_wire_constant when (BITSEL_u8_u1_3064_wire(0) /=  '0') else type_cast_3068_wire_constant;
    -- logger for split-operator MUX_3079_inst flow-through 
    process(IMA76_3080) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3079_inst:flowthrough inputs: " & " BITSEL_u8_u1_3074_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3074_wire) & " type_cast_3076_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3076_wire_constant) & " type_cast_3078_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3078_wire_constant) & " outputs:" & " IMA76_3080= "  & Convert_SLV_To_Hex_String(IMA76_3080));
      --
    end process; 
    -- flow-through select operator MUX_3079_inst
    IMA76_3080 <= type_cast_3076_wire_constant when (BITSEL_u8_u1_3074_wire(0) /=  '0') else type_cast_3078_wire_constant;
    -- logger for split-operator MUX_3089_inst flow-through 
    process(IMA77_3090) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3089_inst:flowthrough inputs: " & " BITSEL_u8_u1_3084_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3084_wire) & " type_cast_3086_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3086_wire_constant) & " type_cast_3088_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3088_wire_constant) & " outputs:" & " IMA77_3090= "  & Convert_SLV_To_Hex_String(IMA77_3090));
      --
    end process; 
    -- flow-through select operator MUX_3089_inst
    IMA77_3090 <= type_cast_3086_wire_constant when (BITSEL_u8_u1_3084_wire(0) /=  '0') else type_cast_3088_wire_constant;
    -- logger for split-operator MUX_3099_inst flow-through 
    process(IMA78_3100) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3099_inst:flowthrough inputs: " & " BITSEL_u8_u1_3094_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3094_wire) & " type_cast_3096_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3096_wire_constant) & " type_cast_3098_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3098_wire_constant) & " outputs:" & " IMA78_3100= "  & Convert_SLV_To_Hex_String(IMA78_3100));
      --
    end process; 
    -- flow-through select operator MUX_3099_inst
    IMA78_3100 <= type_cast_3096_wire_constant when (BITSEL_u8_u1_3094_wire(0) /=  '0') else type_cast_3098_wire_constant;
    -- logger for split-operator MUX_3109_inst flow-through 
    process(IMA79_3110) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3109_inst:flowthrough inputs: " & " BITSEL_u8_u1_3104_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3104_wire) & " type_cast_3106_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3106_wire_constant) & " type_cast_3108_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3108_wire_constant) & " outputs:" & " IMA79_3110= "  & Convert_SLV_To_Hex_String(IMA79_3110));
      --
    end process; 
    -- flow-through select operator MUX_3109_inst
    IMA79_3110 <= type_cast_3106_wire_constant when (BITSEL_u8_u1_3104_wire(0) /=  '0') else type_cast_3108_wire_constant;
    -- logger for split-operator MUX_3119_inst flow-through 
    process(IMA80_3120) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3119_inst:flowthrough inputs: " & " BITSEL_u8_u1_3114_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3114_wire) & " type_cast_3116_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3116_wire_constant) & " type_cast_3118_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3118_wire_constant) & " outputs:" & " IMA80_3120= "  & Convert_SLV_To_Hex_String(IMA80_3120));
      --
    end process; 
    -- flow-through select operator MUX_3119_inst
    IMA80_3120 <= type_cast_3116_wire_constant when (BITSEL_u8_u1_3114_wire(0) /=  '0') else type_cast_3118_wire_constant;
    -- logger for split-operator MUX_3129_inst flow-through 
    process(IMA81_3130) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3129_inst:flowthrough inputs: " & " BITSEL_u8_u1_3124_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3124_wire) & " type_cast_3126_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3126_wire_constant) & " type_cast_3128_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3128_wire_constant) & " outputs:" & " IMA81_3130= "  & Convert_SLV_To_Hex_String(IMA81_3130));
      --
    end process; 
    -- flow-through select operator MUX_3129_inst
    IMA81_3130 <= type_cast_3126_wire_constant when (BITSEL_u8_u1_3124_wire(0) /=  '0') else type_cast_3128_wire_constant;
    -- logger for split-operator MUX_3139_inst flow-through 
    process(IMA82_3140) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3139_inst:flowthrough inputs: " & " BITSEL_u8_u1_3134_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3134_wire) & " type_cast_3136_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3136_wire_constant) & " type_cast_3138_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3138_wire_constant) & " outputs:" & " IMA82_3140= "  & Convert_SLV_To_Hex_String(IMA82_3140));
      --
    end process; 
    -- flow-through select operator MUX_3139_inst
    IMA82_3140 <= type_cast_3136_wire_constant when (BITSEL_u8_u1_3134_wire(0) /=  '0') else type_cast_3138_wire_constant;
    -- logger for split-operator MUX_3149_inst flow-through 
    process(IMA83_3150) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3149_inst:flowthrough inputs: " & " BITSEL_u8_u1_3144_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3144_wire) & " type_cast_3146_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3146_wire_constant) & " type_cast_3148_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3148_wire_constant) & " outputs:" & " IMA83_3150= "  & Convert_SLV_To_Hex_String(IMA83_3150));
      --
    end process; 
    -- flow-through select operator MUX_3149_inst
    IMA83_3150 <= type_cast_3146_wire_constant when (BITSEL_u8_u1_3144_wire(0) /=  '0') else type_cast_3148_wire_constant;
    -- logger for split-operator MUX_3159_inst flow-through 
    process(IMA84_3160) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3159_inst:flowthrough inputs: " & " BITSEL_u8_u1_3154_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3154_wire) & " type_cast_3156_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3156_wire_constant) & " type_cast_3158_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3158_wire_constant) & " outputs:" & " IMA84_3160= "  & Convert_SLV_To_Hex_String(IMA84_3160));
      --
    end process; 
    -- flow-through select operator MUX_3159_inst
    IMA84_3160 <= type_cast_3156_wire_constant when (BITSEL_u8_u1_3154_wire(0) /=  '0') else type_cast_3158_wire_constant;
    -- logger for split-operator MUX_3169_inst flow-through 
    process(IMA85_3170) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3169_inst:flowthrough inputs: " & " BITSEL_u8_u1_3164_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3164_wire) & " type_cast_3166_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3166_wire_constant) & " type_cast_3168_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3168_wire_constant) & " outputs:" & " IMA85_3170= "  & Convert_SLV_To_Hex_String(IMA85_3170));
      --
    end process; 
    -- flow-through select operator MUX_3169_inst
    IMA85_3170 <= type_cast_3166_wire_constant when (BITSEL_u8_u1_3164_wire(0) /=  '0') else type_cast_3168_wire_constant;
    -- logger for split-operator MUX_3179_inst flow-through 
    process(IMA86_3180) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3179_inst:flowthrough inputs: " & " BITSEL_u8_u1_3174_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3174_wire) & " type_cast_3176_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3176_wire_constant) & " type_cast_3178_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3178_wire_constant) & " outputs:" & " IMA86_3180= "  & Convert_SLV_To_Hex_String(IMA86_3180));
      --
    end process; 
    -- flow-through select operator MUX_3179_inst
    IMA86_3180 <= type_cast_3176_wire_constant when (BITSEL_u8_u1_3174_wire(0) /=  '0') else type_cast_3178_wire_constant;
    -- logger for split-operator MUX_3189_inst flow-through 
    process(IMA87_3190) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3189_inst:flowthrough inputs: " & " BITSEL_u8_u1_3184_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3184_wire) & " type_cast_3186_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3186_wire_constant) & " type_cast_3188_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3188_wire_constant) & " outputs:" & " IMA87_3190= "  & Convert_SLV_To_Hex_String(IMA87_3190));
      --
    end process; 
    -- flow-through select operator MUX_3189_inst
    IMA87_3190 <= type_cast_3186_wire_constant when (BITSEL_u8_u1_3184_wire(0) /=  '0') else type_cast_3188_wire_constant;
    -- logger for split-operator MUX_3199_inst flow-through 
    process(IMA88_3200) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3199_inst:flowthrough inputs: " & " BITSEL_u8_u1_3194_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3194_wire) & " type_cast_3196_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3196_wire_constant) & " type_cast_3198_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3198_wire_constant) & " outputs:" & " IMA88_3200= "  & Convert_SLV_To_Hex_String(IMA88_3200));
      --
    end process; 
    -- flow-through select operator MUX_3199_inst
    IMA88_3200 <= type_cast_3196_wire_constant when (BITSEL_u8_u1_3194_wire(0) /=  '0') else type_cast_3198_wire_constant;
    -- logger for split-operator MUX_3209_inst flow-through 
    process(IMA89_3210) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3209_inst:flowthrough inputs: " & " BITSEL_u8_u1_3204_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3204_wire) & " type_cast_3206_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3206_wire_constant) & " type_cast_3208_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3208_wire_constant) & " outputs:" & " IMA89_3210= "  & Convert_SLV_To_Hex_String(IMA89_3210));
      --
    end process; 
    -- flow-through select operator MUX_3209_inst
    IMA89_3210 <= type_cast_3206_wire_constant when (BITSEL_u8_u1_3204_wire(0) /=  '0') else type_cast_3208_wire_constant;
    -- logger for split-operator MUX_3219_inst flow-through 
    process(IMA90_3220) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3219_inst:flowthrough inputs: " & " BITSEL_u8_u1_3214_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3214_wire) & " type_cast_3216_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3216_wire_constant) & " type_cast_3218_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3218_wire_constant) & " outputs:" & " IMA90_3220= "  & Convert_SLV_To_Hex_String(IMA90_3220));
      --
    end process; 
    -- flow-through select operator MUX_3219_inst
    IMA90_3220 <= type_cast_3216_wire_constant when (BITSEL_u8_u1_3214_wire(0) /=  '0') else type_cast_3218_wire_constant;
    -- logger for split-operator MUX_3229_inst flow-through 
    process(IMA91_3230) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3229_inst:flowthrough inputs: " & " BITSEL_u8_u1_3224_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3224_wire) & " type_cast_3226_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3226_wire_constant) & " type_cast_3228_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3228_wire_constant) & " outputs:" & " IMA91_3230= "  & Convert_SLV_To_Hex_String(IMA91_3230));
      --
    end process; 
    -- flow-through select operator MUX_3229_inst
    IMA91_3230 <= type_cast_3226_wire_constant when (BITSEL_u8_u1_3224_wire(0) /=  '0') else type_cast_3228_wire_constant;
    -- logger for split-operator MUX_3239_inst flow-through 
    process(IMA92_3240) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3239_inst:flowthrough inputs: " & " BITSEL_u8_u1_3234_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3234_wire) & " type_cast_3236_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3236_wire_constant) & " type_cast_3238_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3238_wire_constant) & " outputs:" & " IMA92_3240= "  & Convert_SLV_To_Hex_String(IMA92_3240));
      --
    end process; 
    -- flow-through select operator MUX_3239_inst
    IMA92_3240 <= type_cast_3236_wire_constant when (BITSEL_u8_u1_3234_wire(0) /=  '0') else type_cast_3238_wire_constant;
    -- logger for split-operator MUX_3249_inst flow-through 
    process(IMA93_3250) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3249_inst:flowthrough inputs: " & " BITSEL_u8_u1_3244_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3244_wire) & " type_cast_3246_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3246_wire_constant) & " type_cast_3248_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3248_wire_constant) & " outputs:" & " IMA93_3250= "  & Convert_SLV_To_Hex_String(IMA93_3250));
      --
    end process; 
    -- flow-through select operator MUX_3249_inst
    IMA93_3250 <= type_cast_3246_wire_constant when (BITSEL_u8_u1_3244_wire(0) /=  '0') else type_cast_3248_wire_constant;
    -- logger for split-operator MUX_3259_inst flow-through 
    process(IMA94_3260) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3259_inst:flowthrough inputs: " & " BITSEL_u8_u1_3254_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3254_wire) & " type_cast_3256_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3256_wire_constant) & " type_cast_3258_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3258_wire_constant) & " outputs:" & " IMA94_3260= "  & Convert_SLV_To_Hex_String(IMA94_3260));
      --
    end process; 
    -- flow-through select operator MUX_3259_inst
    IMA94_3260 <= type_cast_3256_wire_constant when (BITSEL_u8_u1_3254_wire(0) /=  '0') else type_cast_3258_wire_constant;
    -- logger for split-operator MUX_3269_inst flow-through 
    process(IMA95_3270) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3269_inst:flowthrough inputs: " & " BITSEL_u8_u1_3264_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3264_wire) & " type_cast_3266_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3266_wire_constant) & " type_cast_3268_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3268_wire_constant) & " outputs:" & " IMA95_3270= "  & Convert_SLV_To_Hex_String(IMA95_3270));
      --
    end process; 
    -- flow-through select operator MUX_3269_inst
    IMA95_3270 <= type_cast_3266_wire_constant when (BITSEL_u8_u1_3264_wire(0) /=  '0') else type_cast_3268_wire_constant;
    -- logger for split-operator MUX_3279_inst flow-through 
    process(IMA96_3280) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3279_inst:flowthrough inputs: " & " BITSEL_u8_u1_3274_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3274_wire) & " type_cast_3276_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3276_wire_constant) & " type_cast_3278_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3278_wire_constant) & " outputs:" & " IMA96_3280= "  & Convert_SLV_To_Hex_String(IMA96_3280));
      --
    end process; 
    -- flow-through select operator MUX_3279_inst
    IMA96_3280 <= type_cast_3276_wire_constant when (BITSEL_u8_u1_3274_wire(0) /=  '0') else type_cast_3278_wire_constant;
    -- logger for split-operator MUX_3289_inst flow-through 
    process(IMA97_3290) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3289_inst:flowthrough inputs: " & " BITSEL_u8_u1_3284_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3284_wire) & " type_cast_3286_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3286_wire_constant) & " type_cast_3288_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3288_wire_constant) & " outputs:" & " IMA97_3290= "  & Convert_SLV_To_Hex_String(IMA97_3290));
      --
    end process; 
    -- flow-through select operator MUX_3289_inst
    IMA97_3290 <= type_cast_3286_wire_constant when (BITSEL_u8_u1_3284_wire(0) /=  '0') else type_cast_3288_wire_constant;
    -- logger for split-operator MUX_3299_inst flow-through 
    process(IMA98_3300) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3299_inst:flowthrough inputs: " & " BITSEL_u8_u1_3294_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3294_wire) & " type_cast_3296_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3296_wire_constant) & " type_cast_3298_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3298_wire_constant) & " outputs:" & " IMA98_3300= "  & Convert_SLV_To_Hex_String(IMA98_3300));
      --
    end process; 
    -- flow-through select operator MUX_3299_inst
    IMA98_3300 <= type_cast_3296_wire_constant when (BITSEL_u8_u1_3294_wire(0) /=  '0') else type_cast_3298_wire_constant;
    -- logger for split-operator MUX_3309_inst flow-through 
    process(IMA99_3310) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3309_inst:flowthrough inputs: " & " BITSEL_u8_u1_3304_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3304_wire) & " type_cast_3306_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3306_wire_constant) & " type_cast_3308_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3308_wire_constant) & " outputs:" & " IMA99_3310= "  & Convert_SLV_To_Hex_String(IMA99_3310));
      --
    end process; 
    -- flow-through select operator MUX_3309_inst
    IMA99_3310 <= type_cast_3306_wire_constant when (BITSEL_u8_u1_3304_wire(0) /=  '0') else type_cast_3308_wire_constant;
    -- logger for split-operator MUX_3319_inst flow-through 
    process(IMA100_3320) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3319_inst:flowthrough inputs: " & " BITSEL_u8_u1_3314_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3314_wire) & " type_cast_3316_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3316_wire_constant) & " type_cast_3318_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3318_wire_constant) & " outputs:" & " IMA100_3320= "  & Convert_SLV_To_Hex_String(IMA100_3320));
      --
    end process; 
    -- flow-through select operator MUX_3319_inst
    IMA100_3320 <= type_cast_3316_wire_constant when (BITSEL_u8_u1_3314_wire(0) /=  '0') else type_cast_3318_wire_constant;
    -- logger for split-operator MUX_3329_inst flow-through 
    process(IMA101_3330) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3329_inst:flowthrough inputs: " & " BITSEL_u8_u1_3324_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3324_wire) & " type_cast_3326_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3326_wire_constant) & " type_cast_3328_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3328_wire_constant) & " outputs:" & " IMA101_3330= "  & Convert_SLV_To_Hex_String(IMA101_3330));
      --
    end process; 
    -- flow-through select operator MUX_3329_inst
    IMA101_3330 <= type_cast_3326_wire_constant when (BITSEL_u8_u1_3324_wire(0) /=  '0') else type_cast_3328_wire_constant;
    -- logger for split-operator MUX_3339_inst flow-through 
    process(IMA102_3340) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3339_inst:flowthrough inputs: " & " BITSEL_u8_u1_3334_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3334_wire) & " type_cast_3336_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3336_wire_constant) & " type_cast_3338_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3338_wire_constant) & " outputs:" & " IMA102_3340= "  & Convert_SLV_To_Hex_String(IMA102_3340));
      --
    end process; 
    -- flow-through select operator MUX_3339_inst
    IMA102_3340 <= type_cast_3336_wire_constant when (BITSEL_u8_u1_3334_wire(0) /=  '0') else type_cast_3338_wire_constant;
    -- logger for split-operator MUX_3349_inst flow-through 
    process(IMA103_3350) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3349_inst:flowthrough inputs: " & " BITSEL_u8_u1_3344_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3344_wire) & " type_cast_3346_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3346_wire_constant) & " type_cast_3348_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3348_wire_constant) & " outputs:" & " IMA103_3350= "  & Convert_SLV_To_Hex_String(IMA103_3350));
      --
    end process; 
    -- flow-through select operator MUX_3349_inst
    IMA103_3350 <= type_cast_3346_wire_constant when (BITSEL_u8_u1_3344_wire(0) /=  '0') else type_cast_3348_wire_constant;
    -- logger for split-operator MUX_3359_inst flow-through 
    process(IMA104_3360) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3359_inst:flowthrough inputs: " & " BITSEL_u8_u1_3354_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3354_wire) & " type_cast_3356_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3356_wire_constant) & " type_cast_3358_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3358_wire_constant) & " outputs:" & " IMA104_3360= "  & Convert_SLV_To_Hex_String(IMA104_3360));
      --
    end process; 
    -- flow-through select operator MUX_3359_inst
    IMA104_3360 <= type_cast_3356_wire_constant when (BITSEL_u8_u1_3354_wire(0) /=  '0') else type_cast_3358_wire_constant;
    -- logger for split-operator MUX_3369_inst flow-through 
    process(IMA105_3370) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3369_inst:flowthrough inputs: " & " BITSEL_u8_u1_3364_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3364_wire) & " type_cast_3366_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3366_wire_constant) & " type_cast_3368_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3368_wire_constant) & " outputs:" & " IMA105_3370= "  & Convert_SLV_To_Hex_String(IMA105_3370));
      --
    end process; 
    -- flow-through select operator MUX_3369_inst
    IMA105_3370 <= type_cast_3366_wire_constant when (BITSEL_u8_u1_3364_wire(0) /=  '0') else type_cast_3368_wire_constant;
    -- logger for split-operator MUX_3379_inst flow-through 
    process(IMA106_3380) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3379_inst:flowthrough inputs: " & " BITSEL_u8_u1_3374_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3374_wire) & " type_cast_3376_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3376_wire_constant) & " type_cast_3378_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3378_wire_constant) & " outputs:" & " IMA106_3380= "  & Convert_SLV_To_Hex_String(IMA106_3380));
      --
    end process; 
    -- flow-through select operator MUX_3379_inst
    IMA106_3380 <= type_cast_3376_wire_constant when (BITSEL_u8_u1_3374_wire(0) /=  '0') else type_cast_3378_wire_constant;
    -- logger for split-operator MUX_3389_inst flow-through 
    process(IMA107_3390) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3389_inst:flowthrough inputs: " & " BITSEL_u8_u1_3384_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3384_wire) & " type_cast_3386_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3386_wire_constant) & " type_cast_3388_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3388_wire_constant) & " outputs:" & " IMA107_3390= "  & Convert_SLV_To_Hex_String(IMA107_3390));
      --
    end process; 
    -- flow-through select operator MUX_3389_inst
    IMA107_3390 <= type_cast_3386_wire_constant when (BITSEL_u8_u1_3384_wire(0) /=  '0') else type_cast_3388_wire_constant;
    -- logger for split-operator MUX_3399_inst flow-through 
    process(IMA108_3400) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3399_inst:flowthrough inputs: " & " BITSEL_u8_u1_3394_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3394_wire) & " type_cast_3396_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3396_wire_constant) & " type_cast_3398_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3398_wire_constant) & " outputs:" & " IMA108_3400= "  & Convert_SLV_To_Hex_String(IMA108_3400));
      --
    end process; 
    -- flow-through select operator MUX_3399_inst
    IMA108_3400 <= type_cast_3396_wire_constant when (BITSEL_u8_u1_3394_wire(0) /=  '0') else type_cast_3398_wire_constant;
    -- logger for split-operator MUX_3409_inst flow-through 
    process(IMA109_3410) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3409_inst:flowthrough inputs: " & " BITSEL_u8_u1_3404_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3404_wire) & " type_cast_3406_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3406_wire_constant) & " type_cast_3408_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3408_wire_constant) & " outputs:" & " IMA109_3410= "  & Convert_SLV_To_Hex_String(IMA109_3410));
      --
    end process; 
    -- flow-through select operator MUX_3409_inst
    IMA109_3410 <= type_cast_3406_wire_constant when (BITSEL_u8_u1_3404_wire(0) /=  '0') else type_cast_3408_wire_constant;
    -- logger for split-operator MUX_3419_inst flow-through 
    process(IMA110_3420) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3419_inst:flowthrough inputs: " & " BITSEL_u8_u1_3414_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3414_wire) & " type_cast_3416_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3416_wire_constant) & " type_cast_3418_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3418_wire_constant) & " outputs:" & " IMA110_3420= "  & Convert_SLV_To_Hex_String(IMA110_3420));
      --
    end process; 
    -- flow-through select operator MUX_3419_inst
    IMA110_3420 <= type_cast_3416_wire_constant when (BITSEL_u8_u1_3414_wire(0) /=  '0') else type_cast_3418_wire_constant;
    -- logger for split-operator MUX_3429_inst flow-through 
    process(IMA111_3430) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3429_inst:flowthrough inputs: " & " BITSEL_u8_u1_3424_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3424_wire) & " type_cast_3426_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3426_wire_constant) & " type_cast_3428_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3428_wire_constant) & " outputs:" & " IMA111_3430= "  & Convert_SLV_To_Hex_String(IMA111_3430));
      --
    end process; 
    -- flow-through select operator MUX_3429_inst
    IMA111_3430 <= type_cast_3426_wire_constant when (BITSEL_u8_u1_3424_wire(0) /=  '0') else type_cast_3428_wire_constant;
    -- logger for split-operator MUX_3439_inst flow-through 
    process(IMA112_3440) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3439_inst:flowthrough inputs: " & " BITSEL_u8_u1_3434_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3434_wire) & " type_cast_3436_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3436_wire_constant) & " type_cast_3438_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3438_wire_constant) & " outputs:" & " IMA112_3440= "  & Convert_SLV_To_Hex_String(IMA112_3440));
      --
    end process; 
    -- flow-through select operator MUX_3439_inst
    IMA112_3440 <= type_cast_3436_wire_constant when (BITSEL_u8_u1_3434_wire(0) /=  '0') else type_cast_3438_wire_constant;
    -- logger for split-operator MUX_3449_inst flow-through 
    process(IMA113_3450) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3449_inst:flowthrough inputs: " & " BITSEL_u8_u1_3444_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3444_wire) & " type_cast_3446_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3446_wire_constant) & " type_cast_3448_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3448_wire_constant) & " outputs:" & " IMA113_3450= "  & Convert_SLV_To_Hex_String(IMA113_3450));
      --
    end process; 
    -- flow-through select operator MUX_3449_inst
    IMA113_3450 <= type_cast_3446_wire_constant when (BITSEL_u8_u1_3444_wire(0) /=  '0') else type_cast_3448_wire_constant;
    -- logger for split-operator MUX_3459_inst flow-through 
    process(IMA114_3460) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3459_inst:flowthrough inputs: " & " BITSEL_u8_u1_3454_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3454_wire) & " type_cast_3456_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3456_wire_constant) & " type_cast_3458_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3458_wire_constant) & " outputs:" & " IMA114_3460= "  & Convert_SLV_To_Hex_String(IMA114_3460));
      --
    end process; 
    -- flow-through select operator MUX_3459_inst
    IMA114_3460 <= type_cast_3456_wire_constant when (BITSEL_u8_u1_3454_wire(0) /=  '0') else type_cast_3458_wire_constant;
    -- logger for split-operator MUX_3469_inst flow-through 
    process(IMA115_3470) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3469_inst:flowthrough inputs: " & " BITSEL_u8_u1_3464_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3464_wire) & " type_cast_3466_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3466_wire_constant) & " type_cast_3468_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3468_wire_constant) & " outputs:" & " IMA115_3470= "  & Convert_SLV_To_Hex_String(IMA115_3470));
      --
    end process; 
    -- flow-through select operator MUX_3469_inst
    IMA115_3470 <= type_cast_3466_wire_constant when (BITSEL_u8_u1_3464_wire(0) /=  '0') else type_cast_3468_wire_constant;
    -- logger for split-operator MUX_3479_inst flow-through 
    process(IMA116_3480) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3479_inst:flowthrough inputs: " & " BITSEL_u8_u1_3474_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3474_wire) & " type_cast_3476_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3476_wire_constant) & " type_cast_3478_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3478_wire_constant) & " outputs:" & " IMA116_3480= "  & Convert_SLV_To_Hex_String(IMA116_3480));
      --
    end process; 
    -- flow-through select operator MUX_3479_inst
    IMA116_3480 <= type_cast_3476_wire_constant when (BITSEL_u8_u1_3474_wire(0) /=  '0') else type_cast_3478_wire_constant;
    -- logger for split-operator MUX_3489_inst flow-through 
    process(IMA117_3490) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3489_inst:flowthrough inputs: " & " BITSEL_u8_u1_3484_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3484_wire) & " type_cast_3486_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3486_wire_constant) & " type_cast_3488_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3488_wire_constant) & " outputs:" & " IMA117_3490= "  & Convert_SLV_To_Hex_String(IMA117_3490));
      --
    end process; 
    -- flow-through select operator MUX_3489_inst
    IMA117_3490 <= type_cast_3486_wire_constant when (BITSEL_u8_u1_3484_wire(0) /=  '0') else type_cast_3488_wire_constant;
    -- logger for split-operator MUX_3499_inst flow-through 
    process(IMA118_3500) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3499_inst:flowthrough inputs: " & " BITSEL_u8_u1_3494_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3494_wire) & " type_cast_3496_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3496_wire_constant) & " type_cast_3498_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3498_wire_constant) & " outputs:" & " IMA118_3500= "  & Convert_SLV_To_Hex_String(IMA118_3500));
      --
    end process; 
    -- flow-through select operator MUX_3499_inst
    IMA118_3500 <= type_cast_3496_wire_constant when (BITSEL_u8_u1_3494_wire(0) /=  '0') else type_cast_3498_wire_constant;
    -- logger for split-operator MUX_3509_inst flow-through 
    process(IMA119_3510) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3509_inst:flowthrough inputs: " & " BITSEL_u8_u1_3504_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3504_wire) & " type_cast_3506_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3506_wire_constant) & " type_cast_3508_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3508_wire_constant) & " outputs:" & " IMA119_3510= "  & Convert_SLV_To_Hex_String(IMA119_3510));
      --
    end process; 
    -- flow-through select operator MUX_3509_inst
    IMA119_3510 <= type_cast_3506_wire_constant when (BITSEL_u8_u1_3504_wire(0) /=  '0') else type_cast_3508_wire_constant;
    -- logger for split-operator MUX_3519_inst flow-through 
    process(IMA120_3520) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3519_inst:flowthrough inputs: " & " BITSEL_u8_u1_3514_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3514_wire) & " type_cast_3516_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3516_wire_constant) & " type_cast_3518_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3518_wire_constant) & " outputs:" & " IMA120_3520= "  & Convert_SLV_To_Hex_String(IMA120_3520));
      --
    end process; 
    -- flow-through select operator MUX_3519_inst
    IMA120_3520 <= type_cast_3516_wire_constant when (BITSEL_u8_u1_3514_wire(0) /=  '0') else type_cast_3518_wire_constant;
    -- logger for split-operator MUX_3529_inst flow-through 
    process(IMA121_3530) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3529_inst:flowthrough inputs: " & " BITSEL_u8_u1_3524_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3524_wire) & " type_cast_3526_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3526_wire_constant) & " type_cast_3528_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3528_wire_constant) & " outputs:" & " IMA121_3530= "  & Convert_SLV_To_Hex_String(IMA121_3530));
      --
    end process; 
    -- flow-through select operator MUX_3529_inst
    IMA121_3530 <= type_cast_3526_wire_constant when (BITSEL_u8_u1_3524_wire(0) /=  '0') else type_cast_3528_wire_constant;
    -- logger for split-operator MUX_3539_inst flow-through 
    process(IMA122_3540) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3539_inst:flowthrough inputs: " & " BITSEL_u8_u1_3534_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3534_wire) & " type_cast_3536_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3536_wire_constant) & " type_cast_3538_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3538_wire_constant) & " outputs:" & " IMA122_3540= "  & Convert_SLV_To_Hex_String(IMA122_3540));
      --
    end process; 
    -- flow-through select operator MUX_3539_inst
    IMA122_3540 <= type_cast_3536_wire_constant when (BITSEL_u8_u1_3534_wire(0) /=  '0') else type_cast_3538_wire_constant;
    -- logger for split-operator MUX_3549_inst flow-through 
    process(IMA123_3550) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3549_inst:flowthrough inputs: " & " BITSEL_u8_u1_3544_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3544_wire) & " type_cast_3546_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3546_wire_constant) & " type_cast_3548_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3548_wire_constant) & " outputs:" & " IMA123_3550= "  & Convert_SLV_To_Hex_String(IMA123_3550));
      --
    end process; 
    -- flow-through select operator MUX_3549_inst
    IMA123_3550 <= type_cast_3546_wire_constant when (BITSEL_u8_u1_3544_wire(0) /=  '0') else type_cast_3548_wire_constant;
    -- logger for split-operator MUX_3559_inst flow-through 
    process(IMA124_3560) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3559_inst:flowthrough inputs: " & " BITSEL_u8_u1_3554_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3554_wire) & " type_cast_3556_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3556_wire_constant) & " type_cast_3558_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3558_wire_constant) & " outputs:" & " IMA124_3560= "  & Convert_SLV_To_Hex_String(IMA124_3560));
      --
    end process; 
    -- flow-through select operator MUX_3559_inst
    IMA124_3560 <= type_cast_3556_wire_constant when (BITSEL_u8_u1_3554_wire(0) /=  '0') else type_cast_3558_wire_constant;
    -- logger for split-operator MUX_3569_inst flow-through 
    process(IMA125_3570) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3569_inst:flowthrough inputs: " & " BITSEL_u8_u1_3564_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3564_wire) & " type_cast_3566_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3566_wire_constant) & " type_cast_3568_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3568_wire_constant) & " outputs:" & " IMA125_3570= "  & Convert_SLV_To_Hex_String(IMA125_3570));
      --
    end process; 
    -- flow-through select operator MUX_3569_inst
    IMA125_3570 <= type_cast_3566_wire_constant when (BITSEL_u8_u1_3564_wire(0) /=  '0') else type_cast_3568_wire_constant;
    -- logger for split-operator MUX_3579_inst flow-through 
    process(IMA126_3580) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3579_inst:flowthrough inputs: " & " BITSEL_u8_u1_3574_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3574_wire) & " type_cast_3576_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3576_wire_constant) & " type_cast_3578_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3578_wire_constant) & " outputs:" & " IMA126_3580= "  & Convert_SLV_To_Hex_String(IMA126_3580));
      --
    end process; 
    -- flow-through select operator MUX_3579_inst
    IMA126_3580 <= type_cast_3576_wire_constant when (BITSEL_u8_u1_3574_wire(0) /=  '0') else type_cast_3578_wire_constant;
    -- logger for split-operator MUX_3589_inst flow-through 
    process(IMA127_3590) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3589_inst:flowthrough inputs: " & " BITSEL_u8_u1_3584_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3584_wire) & " type_cast_3586_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3586_wire_constant) & " type_cast_3588_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_3588_wire_constant) & " outputs:" & " IMA127_3590= "  & Convert_SLV_To_Hex_String(IMA127_3590));
      --
    end process; 
    -- flow-through select operator MUX_3589_inst
    IMA127_3590 <= type_cast_3586_wire_constant when (BITSEL_u8_u1_3584_wire(0) /=  '0') else type_cast_3588_wire_constant;
    -- logger for split-operator MUX_3597_inst flow-through 
    process(IMB0_3598) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3597_inst:flowthrough inputs: " & " BITSEL_u8_u1_3594_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3594_wire) & " IMA1_2330 = "& Convert_SLV_To_Hex_String(IMA1_2330) & " IMA0_2320 = "& Convert_SLV_To_Hex_String(IMA0_2320) & " outputs:" & " IMB0_3598= "  & Convert_SLV_To_Hex_String(IMB0_3598));
      --
    end process; 
    -- flow-through select operator MUX_3597_inst
    IMB0_3598 <= IMA1_2330 when (BITSEL_u8_u1_3594_wire(0) /=  '0') else IMA0_2320;
    -- logger for split-operator MUX_3605_inst flow-through 
    process(IMB1_3606) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3605_inst:flowthrough inputs: " & " BITSEL_u8_u1_3602_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3602_wire) & " IMA3_2350 = "& Convert_SLV_To_Hex_String(IMA3_2350) & " IMA2_2340 = "& Convert_SLV_To_Hex_String(IMA2_2340) & " outputs:" & " IMB1_3606= "  & Convert_SLV_To_Hex_String(IMB1_3606));
      --
    end process; 
    -- flow-through select operator MUX_3605_inst
    IMB1_3606 <= IMA3_2350 when (BITSEL_u8_u1_3602_wire(0) /=  '0') else IMA2_2340;
    -- logger for split-operator MUX_3613_inst flow-through 
    process(IMB2_3614) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3613_inst:flowthrough inputs: " & " BITSEL_u8_u1_3610_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3610_wire) & " IMA5_2370 = "& Convert_SLV_To_Hex_String(IMA5_2370) & " IMA4_2360 = "& Convert_SLV_To_Hex_String(IMA4_2360) & " outputs:" & " IMB2_3614= "  & Convert_SLV_To_Hex_String(IMB2_3614));
      --
    end process; 
    -- flow-through select operator MUX_3613_inst
    IMB2_3614 <= IMA5_2370 when (BITSEL_u8_u1_3610_wire(0) /=  '0') else IMA4_2360;
    -- logger for split-operator MUX_3621_inst flow-through 
    process(IMB3_3622) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3621_inst:flowthrough inputs: " & " BITSEL_u8_u1_3618_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3618_wire) & " IMA7_2390 = "& Convert_SLV_To_Hex_String(IMA7_2390) & " IMA6_2380 = "& Convert_SLV_To_Hex_String(IMA6_2380) & " outputs:" & " IMB3_3622= "  & Convert_SLV_To_Hex_String(IMB3_3622));
      --
    end process; 
    -- flow-through select operator MUX_3621_inst
    IMB3_3622 <= IMA7_2390 when (BITSEL_u8_u1_3618_wire(0) /=  '0') else IMA6_2380;
    -- logger for split-operator MUX_3629_inst flow-through 
    process(IMB4_3630) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3629_inst:flowthrough inputs: " & " BITSEL_u8_u1_3626_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3626_wire) & " IMA9_2410 = "& Convert_SLV_To_Hex_String(IMA9_2410) & " IMA8_2400 = "& Convert_SLV_To_Hex_String(IMA8_2400) & " outputs:" & " IMB4_3630= "  & Convert_SLV_To_Hex_String(IMB4_3630));
      --
    end process; 
    -- flow-through select operator MUX_3629_inst
    IMB4_3630 <= IMA9_2410 when (BITSEL_u8_u1_3626_wire(0) /=  '0') else IMA8_2400;
    -- logger for split-operator MUX_3637_inst flow-through 
    process(IMB5_3638) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3637_inst:flowthrough inputs: " & " BITSEL_u8_u1_3634_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3634_wire) & " IMA11_2430 = "& Convert_SLV_To_Hex_String(IMA11_2430) & " IMA10_2420 = "& Convert_SLV_To_Hex_String(IMA10_2420) & " outputs:" & " IMB5_3638= "  & Convert_SLV_To_Hex_String(IMB5_3638));
      --
    end process; 
    -- flow-through select operator MUX_3637_inst
    IMB5_3638 <= IMA11_2430 when (BITSEL_u8_u1_3634_wire(0) /=  '0') else IMA10_2420;
    -- logger for split-operator MUX_3645_inst flow-through 
    process(IMB6_3646) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3645_inst:flowthrough inputs: " & " BITSEL_u8_u1_3642_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3642_wire) & " IMA13_2450 = "& Convert_SLV_To_Hex_String(IMA13_2450) & " IMA12_2440 = "& Convert_SLV_To_Hex_String(IMA12_2440) & " outputs:" & " IMB6_3646= "  & Convert_SLV_To_Hex_String(IMB6_3646));
      --
    end process; 
    -- flow-through select operator MUX_3645_inst
    IMB6_3646 <= IMA13_2450 when (BITSEL_u8_u1_3642_wire(0) /=  '0') else IMA12_2440;
    -- logger for split-operator MUX_3653_inst flow-through 
    process(IMB7_3654) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3653_inst:flowthrough inputs: " & " BITSEL_u8_u1_3650_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3650_wire) & " IMA15_2470 = "& Convert_SLV_To_Hex_String(IMA15_2470) & " IMA14_2460 = "& Convert_SLV_To_Hex_String(IMA14_2460) & " outputs:" & " IMB7_3654= "  & Convert_SLV_To_Hex_String(IMB7_3654));
      --
    end process; 
    -- flow-through select operator MUX_3653_inst
    IMB7_3654 <= IMA15_2470 when (BITSEL_u8_u1_3650_wire(0) /=  '0') else IMA14_2460;
    -- logger for split-operator MUX_3661_inst flow-through 
    process(IMB8_3662) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3661_inst:flowthrough inputs: " & " BITSEL_u8_u1_3658_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3658_wire) & " IMA17_2490 = "& Convert_SLV_To_Hex_String(IMA17_2490) & " IMA16_2480 = "& Convert_SLV_To_Hex_String(IMA16_2480) & " outputs:" & " IMB8_3662= "  & Convert_SLV_To_Hex_String(IMB8_3662));
      --
    end process; 
    -- flow-through select operator MUX_3661_inst
    IMB8_3662 <= IMA17_2490 when (BITSEL_u8_u1_3658_wire(0) /=  '0') else IMA16_2480;
    -- logger for split-operator MUX_3669_inst flow-through 
    process(IMB9_3670) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3669_inst:flowthrough inputs: " & " BITSEL_u8_u1_3666_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3666_wire) & " IMA19_2510 = "& Convert_SLV_To_Hex_String(IMA19_2510) & " IMA18_2500 = "& Convert_SLV_To_Hex_String(IMA18_2500) & " outputs:" & " IMB9_3670= "  & Convert_SLV_To_Hex_String(IMB9_3670));
      --
    end process; 
    -- flow-through select operator MUX_3669_inst
    IMB9_3670 <= IMA19_2510 when (BITSEL_u8_u1_3666_wire(0) /=  '0') else IMA18_2500;
    -- logger for split-operator MUX_3677_inst flow-through 
    process(IMB10_3678) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3677_inst:flowthrough inputs: " & " BITSEL_u8_u1_3674_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3674_wire) & " IMA21_2530 = "& Convert_SLV_To_Hex_String(IMA21_2530) & " IMA20_2520 = "& Convert_SLV_To_Hex_String(IMA20_2520) & " outputs:" & " IMB10_3678= "  & Convert_SLV_To_Hex_String(IMB10_3678));
      --
    end process; 
    -- flow-through select operator MUX_3677_inst
    IMB10_3678 <= IMA21_2530 when (BITSEL_u8_u1_3674_wire(0) /=  '0') else IMA20_2520;
    -- logger for split-operator MUX_3685_inst flow-through 
    process(IMB11_3686) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3685_inst:flowthrough inputs: " & " BITSEL_u8_u1_3682_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3682_wire) & " IMA23_2550 = "& Convert_SLV_To_Hex_String(IMA23_2550) & " IMA22_2540 = "& Convert_SLV_To_Hex_String(IMA22_2540) & " outputs:" & " IMB11_3686= "  & Convert_SLV_To_Hex_String(IMB11_3686));
      --
    end process; 
    -- flow-through select operator MUX_3685_inst
    IMB11_3686 <= IMA23_2550 when (BITSEL_u8_u1_3682_wire(0) /=  '0') else IMA22_2540;
    -- logger for split-operator MUX_3693_inst flow-through 
    process(IMB12_3694) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3693_inst:flowthrough inputs: " & " BITSEL_u8_u1_3690_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3690_wire) & " IMA25_2570 = "& Convert_SLV_To_Hex_String(IMA25_2570) & " IMA24_2560 = "& Convert_SLV_To_Hex_String(IMA24_2560) & " outputs:" & " IMB12_3694= "  & Convert_SLV_To_Hex_String(IMB12_3694));
      --
    end process; 
    -- flow-through select operator MUX_3693_inst
    IMB12_3694 <= IMA25_2570 when (BITSEL_u8_u1_3690_wire(0) /=  '0') else IMA24_2560;
    -- logger for split-operator MUX_3701_inst flow-through 
    process(IMB13_3702) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3701_inst:flowthrough inputs: " & " BITSEL_u8_u1_3698_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3698_wire) & " IMA27_2590 = "& Convert_SLV_To_Hex_String(IMA27_2590) & " IMA26_2580 = "& Convert_SLV_To_Hex_String(IMA26_2580) & " outputs:" & " IMB13_3702= "  & Convert_SLV_To_Hex_String(IMB13_3702));
      --
    end process; 
    -- flow-through select operator MUX_3701_inst
    IMB13_3702 <= IMA27_2590 when (BITSEL_u8_u1_3698_wire(0) /=  '0') else IMA26_2580;
    -- logger for split-operator MUX_3709_inst flow-through 
    process(IMB14_3710) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3709_inst:flowthrough inputs: " & " BITSEL_u8_u1_3706_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3706_wire) & " IMA29_2610 = "& Convert_SLV_To_Hex_String(IMA29_2610) & " IMA28_2600 = "& Convert_SLV_To_Hex_String(IMA28_2600) & " outputs:" & " IMB14_3710= "  & Convert_SLV_To_Hex_String(IMB14_3710));
      --
    end process; 
    -- flow-through select operator MUX_3709_inst
    IMB14_3710 <= IMA29_2610 when (BITSEL_u8_u1_3706_wire(0) /=  '0') else IMA28_2600;
    -- logger for split-operator MUX_3717_inst flow-through 
    process(IMB15_3718) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3717_inst:flowthrough inputs: " & " BITSEL_u8_u1_3714_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3714_wire) & " IMA31_2630 = "& Convert_SLV_To_Hex_String(IMA31_2630) & " IMA30_2620 = "& Convert_SLV_To_Hex_String(IMA30_2620) & " outputs:" & " IMB15_3718= "  & Convert_SLV_To_Hex_String(IMB15_3718));
      --
    end process; 
    -- flow-through select operator MUX_3717_inst
    IMB15_3718 <= IMA31_2630 when (BITSEL_u8_u1_3714_wire(0) /=  '0') else IMA30_2620;
    -- logger for split-operator MUX_3725_inst flow-through 
    process(IMB16_3726) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3725_inst:flowthrough inputs: " & " BITSEL_u8_u1_3722_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3722_wire) & " IMA33_2650 = "& Convert_SLV_To_Hex_String(IMA33_2650) & " IMA32_2640 = "& Convert_SLV_To_Hex_String(IMA32_2640) & " outputs:" & " IMB16_3726= "  & Convert_SLV_To_Hex_String(IMB16_3726));
      --
    end process; 
    -- flow-through select operator MUX_3725_inst
    IMB16_3726 <= IMA33_2650 when (BITSEL_u8_u1_3722_wire(0) /=  '0') else IMA32_2640;
    -- logger for split-operator MUX_3733_inst flow-through 
    process(IMB17_3734) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3733_inst:flowthrough inputs: " & " BITSEL_u8_u1_3730_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3730_wire) & " IMA35_2670 = "& Convert_SLV_To_Hex_String(IMA35_2670) & " IMA34_2660 = "& Convert_SLV_To_Hex_String(IMA34_2660) & " outputs:" & " IMB17_3734= "  & Convert_SLV_To_Hex_String(IMB17_3734));
      --
    end process; 
    -- flow-through select operator MUX_3733_inst
    IMB17_3734 <= IMA35_2670 when (BITSEL_u8_u1_3730_wire(0) /=  '0') else IMA34_2660;
    -- logger for split-operator MUX_3741_inst flow-through 
    process(IMB18_3742) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3741_inst:flowthrough inputs: " & " BITSEL_u8_u1_3738_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3738_wire) & " IMA37_2690 = "& Convert_SLV_To_Hex_String(IMA37_2690) & " IMA36_2680 = "& Convert_SLV_To_Hex_String(IMA36_2680) & " outputs:" & " IMB18_3742= "  & Convert_SLV_To_Hex_String(IMB18_3742));
      --
    end process; 
    -- flow-through select operator MUX_3741_inst
    IMB18_3742 <= IMA37_2690 when (BITSEL_u8_u1_3738_wire(0) /=  '0') else IMA36_2680;
    -- logger for split-operator MUX_3749_inst flow-through 
    process(IMB19_3750) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3749_inst:flowthrough inputs: " & " BITSEL_u8_u1_3746_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3746_wire) & " IMA39_2710 = "& Convert_SLV_To_Hex_String(IMA39_2710) & " IMA38_2700 = "& Convert_SLV_To_Hex_String(IMA38_2700) & " outputs:" & " IMB19_3750= "  & Convert_SLV_To_Hex_String(IMB19_3750));
      --
    end process; 
    -- flow-through select operator MUX_3749_inst
    IMB19_3750 <= IMA39_2710 when (BITSEL_u8_u1_3746_wire(0) /=  '0') else IMA38_2700;
    -- logger for split-operator MUX_3757_inst flow-through 
    process(IMB20_3758) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3757_inst:flowthrough inputs: " & " BITSEL_u8_u1_3754_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3754_wire) & " IMA41_2730 = "& Convert_SLV_To_Hex_String(IMA41_2730) & " IMA40_2720 = "& Convert_SLV_To_Hex_String(IMA40_2720) & " outputs:" & " IMB20_3758= "  & Convert_SLV_To_Hex_String(IMB20_3758));
      --
    end process; 
    -- flow-through select operator MUX_3757_inst
    IMB20_3758 <= IMA41_2730 when (BITSEL_u8_u1_3754_wire(0) /=  '0') else IMA40_2720;
    -- logger for split-operator MUX_3765_inst flow-through 
    process(IMB21_3766) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3765_inst:flowthrough inputs: " & " BITSEL_u8_u1_3762_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3762_wire) & " IMA43_2750 = "& Convert_SLV_To_Hex_String(IMA43_2750) & " IMA42_2740 = "& Convert_SLV_To_Hex_String(IMA42_2740) & " outputs:" & " IMB21_3766= "  & Convert_SLV_To_Hex_String(IMB21_3766));
      --
    end process; 
    -- flow-through select operator MUX_3765_inst
    IMB21_3766 <= IMA43_2750 when (BITSEL_u8_u1_3762_wire(0) /=  '0') else IMA42_2740;
    -- logger for split-operator MUX_3773_inst flow-through 
    process(IMB22_3774) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3773_inst:flowthrough inputs: " & " BITSEL_u8_u1_3770_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3770_wire) & " IMA45_2770 = "& Convert_SLV_To_Hex_String(IMA45_2770) & " IMA44_2760 = "& Convert_SLV_To_Hex_String(IMA44_2760) & " outputs:" & " IMB22_3774= "  & Convert_SLV_To_Hex_String(IMB22_3774));
      --
    end process; 
    -- flow-through select operator MUX_3773_inst
    IMB22_3774 <= IMA45_2770 when (BITSEL_u8_u1_3770_wire(0) /=  '0') else IMA44_2760;
    -- logger for split-operator MUX_3781_inst flow-through 
    process(IMB23_3782) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3781_inst:flowthrough inputs: " & " BITSEL_u8_u1_3778_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3778_wire) & " IMA47_2790 = "& Convert_SLV_To_Hex_String(IMA47_2790) & " IMA46_2780 = "& Convert_SLV_To_Hex_String(IMA46_2780) & " outputs:" & " IMB23_3782= "  & Convert_SLV_To_Hex_String(IMB23_3782));
      --
    end process; 
    -- flow-through select operator MUX_3781_inst
    IMB23_3782 <= IMA47_2790 when (BITSEL_u8_u1_3778_wire(0) /=  '0') else IMA46_2780;
    -- logger for split-operator MUX_3789_inst flow-through 
    process(IMB24_3790) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3789_inst:flowthrough inputs: " & " BITSEL_u8_u1_3786_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3786_wire) & " IMA49_2810 = "& Convert_SLV_To_Hex_String(IMA49_2810) & " IMA48_2800 = "& Convert_SLV_To_Hex_String(IMA48_2800) & " outputs:" & " IMB24_3790= "  & Convert_SLV_To_Hex_String(IMB24_3790));
      --
    end process; 
    -- flow-through select operator MUX_3789_inst
    IMB24_3790 <= IMA49_2810 when (BITSEL_u8_u1_3786_wire(0) /=  '0') else IMA48_2800;
    -- logger for split-operator MUX_3797_inst flow-through 
    process(IMB25_3798) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3797_inst:flowthrough inputs: " & " BITSEL_u8_u1_3794_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3794_wire) & " IMA51_2830 = "& Convert_SLV_To_Hex_String(IMA51_2830) & " IMA50_2820 = "& Convert_SLV_To_Hex_String(IMA50_2820) & " outputs:" & " IMB25_3798= "  & Convert_SLV_To_Hex_String(IMB25_3798));
      --
    end process; 
    -- flow-through select operator MUX_3797_inst
    IMB25_3798 <= IMA51_2830 when (BITSEL_u8_u1_3794_wire(0) /=  '0') else IMA50_2820;
    -- logger for split-operator MUX_3805_inst flow-through 
    process(IMB26_3806) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3805_inst:flowthrough inputs: " & " BITSEL_u8_u1_3802_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3802_wire) & " IMA53_2850 = "& Convert_SLV_To_Hex_String(IMA53_2850) & " IMA52_2840 = "& Convert_SLV_To_Hex_String(IMA52_2840) & " outputs:" & " IMB26_3806= "  & Convert_SLV_To_Hex_String(IMB26_3806));
      --
    end process; 
    -- flow-through select operator MUX_3805_inst
    IMB26_3806 <= IMA53_2850 when (BITSEL_u8_u1_3802_wire(0) /=  '0') else IMA52_2840;
    -- logger for split-operator MUX_3813_inst flow-through 
    process(IMB27_3814) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3813_inst:flowthrough inputs: " & " BITSEL_u8_u1_3810_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3810_wire) & " IMA55_2870 = "& Convert_SLV_To_Hex_String(IMA55_2870) & " IMA54_2860 = "& Convert_SLV_To_Hex_String(IMA54_2860) & " outputs:" & " IMB27_3814= "  & Convert_SLV_To_Hex_String(IMB27_3814));
      --
    end process; 
    -- flow-through select operator MUX_3813_inst
    IMB27_3814 <= IMA55_2870 when (BITSEL_u8_u1_3810_wire(0) /=  '0') else IMA54_2860;
    -- logger for split-operator MUX_3821_inst flow-through 
    process(IMB28_3822) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3821_inst:flowthrough inputs: " & " BITSEL_u8_u1_3818_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3818_wire) & " IMA57_2890 = "& Convert_SLV_To_Hex_String(IMA57_2890) & " IMA56_2880 = "& Convert_SLV_To_Hex_String(IMA56_2880) & " outputs:" & " IMB28_3822= "  & Convert_SLV_To_Hex_String(IMB28_3822));
      --
    end process; 
    -- flow-through select operator MUX_3821_inst
    IMB28_3822 <= IMA57_2890 when (BITSEL_u8_u1_3818_wire(0) /=  '0') else IMA56_2880;
    -- logger for split-operator MUX_3829_inst flow-through 
    process(IMB29_3830) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3829_inst:flowthrough inputs: " & " BITSEL_u8_u1_3826_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3826_wire) & " IMA59_2910 = "& Convert_SLV_To_Hex_String(IMA59_2910) & " IMA58_2900 = "& Convert_SLV_To_Hex_String(IMA58_2900) & " outputs:" & " IMB29_3830= "  & Convert_SLV_To_Hex_String(IMB29_3830));
      --
    end process; 
    -- flow-through select operator MUX_3829_inst
    IMB29_3830 <= IMA59_2910 when (BITSEL_u8_u1_3826_wire(0) /=  '0') else IMA58_2900;
    -- logger for split-operator MUX_3837_inst flow-through 
    process(IMB30_3838) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3837_inst:flowthrough inputs: " & " BITSEL_u8_u1_3834_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3834_wire) & " IMA61_2930 = "& Convert_SLV_To_Hex_String(IMA61_2930) & " IMA60_2920 = "& Convert_SLV_To_Hex_String(IMA60_2920) & " outputs:" & " IMB30_3838= "  & Convert_SLV_To_Hex_String(IMB30_3838));
      --
    end process; 
    -- flow-through select operator MUX_3837_inst
    IMB30_3838 <= IMA61_2930 when (BITSEL_u8_u1_3834_wire(0) /=  '0') else IMA60_2920;
    -- logger for split-operator MUX_3845_inst flow-through 
    process(IMB31_3846) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3845_inst:flowthrough inputs: " & " BITSEL_u8_u1_3842_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3842_wire) & " IMA63_2950 = "& Convert_SLV_To_Hex_String(IMA63_2950) & " IMA62_2940 = "& Convert_SLV_To_Hex_String(IMA62_2940) & " outputs:" & " IMB31_3846= "  & Convert_SLV_To_Hex_String(IMB31_3846));
      --
    end process; 
    -- flow-through select operator MUX_3845_inst
    IMB31_3846 <= IMA63_2950 when (BITSEL_u8_u1_3842_wire(0) /=  '0') else IMA62_2940;
    -- logger for split-operator MUX_3853_inst flow-through 
    process(IMB32_3854) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3853_inst:flowthrough inputs: " & " BITSEL_u8_u1_3850_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3850_wire) & " IMA65_2970 = "& Convert_SLV_To_Hex_String(IMA65_2970) & " IMA64_2960 = "& Convert_SLV_To_Hex_String(IMA64_2960) & " outputs:" & " IMB32_3854= "  & Convert_SLV_To_Hex_String(IMB32_3854));
      --
    end process; 
    -- flow-through select operator MUX_3853_inst
    IMB32_3854 <= IMA65_2970 when (BITSEL_u8_u1_3850_wire(0) /=  '0') else IMA64_2960;
    -- logger for split-operator MUX_3861_inst flow-through 
    process(IMB33_3862) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3861_inst:flowthrough inputs: " & " BITSEL_u8_u1_3858_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3858_wire) & " IMA67_2990 = "& Convert_SLV_To_Hex_String(IMA67_2990) & " IMA66_2980 = "& Convert_SLV_To_Hex_String(IMA66_2980) & " outputs:" & " IMB33_3862= "  & Convert_SLV_To_Hex_String(IMB33_3862));
      --
    end process; 
    -- flow-through select operator MUX_3861_inst
    IMB33_3862 <= IMA67_2990 when (BITSEL_u8_u1_3858_wire(0) /=  '0') else IMA66_2980;
    -- logger for split-operator MUX_3869_inst flow-through 
    process(IMB34_3870) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3869_inst:flowthrough inputs: " & " BITSEL_u8_u1_3866_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3866_wire) & " IMA69_3010 = "& Convert_SLV_To_Hex_String(IMA69_3010) & " IMA68_3000 = "& Convert_SLV_To_Hex_String(IMA68_3000) & " outputs:" & " IMB34_3870= "  & Convert_SLV_To_Hex_String(IMB34_3870));
      --
    end process; 
    -- flow-through select operator MUX_3869_inst
    IMB34_3870 <= IMA69_3010 when (BITSEL_u8_u1_3866_wire(0) /=  '0') else IMA68_3000;
    -- logger for split-operator MUX_3877_inst flow-through 
    process(IMB35_3878) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3877_inst:flowthrough inputs: " & " BITSEL_u8_u1_3874_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3874_wire) & " IMA71_3030 = "& Convert_SLV_To_Hex_String(IMA71_3030) & " IMA70_3020 = "& Convert_SLV_To_Hex_String(IMA70_3020) & " outputs:" & " IMB35_3878= "  & Convert_SLV_To_Hex_String(IMB35_3878));
      --
    end process; 
    -- flow-through select operator MUX_3877_inst
    IMB35_3878 <= IMA71_3030 when (BITSEL_u8_u1_3874_wire(0) /=  '0') else IMA70_3020;
    -- logger for split-operator MUX_3885_inst flow-through 
    process(IMB36_3886) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3885_inst:flowthrough inputs: " & " BITSEL_u8_u1_3882_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3882_wire) & " IMA73_3050 = "& Convert_SLV_To_Hex_String(IMA73_3050) & " IMA72_3040 = "& Convert_SLV_To_Hex_String(IMA72_3040) & " outputs:" & " IMB36_3886= "  & Convert_SLV_To_Hex_String(IMB36_3886));
      --
    end process; 
    -- flow-through select operator MUX_3885_inst
    IMB36_3886 <= IMA73_3050 when (BITSEL_u8_u1_3882_wire(0) /=  '0') else IMA72_3040;
    -- logger for split-operator MUX_3893_inst flow-through 
    process(IMB37_3894) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3893_inst:flowthrough inputs: " & " BITSEL_u8_u1_3890_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3890_wire) & " IMA75_3070 = "& Convert_SLV_To_Hex_String(IMA75_3070) & " IMA74_3060 = "& Convert_SLV_To_Hex_String(IMA74_3060) & " outputs:" & " IMB37_3894= "  & Convert_SLV_To_Hex_String(IMB37_3894));
      --
    end process; 
    -- flow-through select operator MUX_3893_inst
    IMB37_3894 <= IMA75_3070 when (BITSEL_u8_u1_3890_wire(0) /=  '0') else IMA74_3060;
    -- logger for split-operator MUX_3901_inst flow-through 
    process(IMB38_3902) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3901_inst:flowthrough inputs: " & " BITSEL_u8_u1_3898_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3898_wire) & " IMA77_3090 = "& Convert_SLV_To_Hex_String(IMA77_3090) & " IMA76_3080 = "& Convert_SLV_To_Hex_String(IMA76_3080) & " outputs:" & " IMB38_3902= "  & Convert_SLV_To_Hex_String(IMB38_3902));
      --
    end process; 
    -- flow-through select operator MUX_3901_inst
    IMB38_3902 <= IMA77_3090 when (BITSEL_u8_u1_3898_wire(0) /=  '0') else IMA76_3080;
    -- logger for split-operator MUX_3909_inst flow-through 
    process(IMB39_3910) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3909_inst:flowthrough inputs: " & " BITSEL_u8_u1_3906_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3906_wire) & " IMA79_3110 = "& Convert_SLV_To_Hex_String(IMA79_3110) & " IMA78_3100 = "& Convert_SLV_To_Hex_String(IMA78_3100) & " outputs:" & " IMB39_3910= "  & Convert_SLV_To_Hex_String(IMB39_3910));
      --
    end process; 
    -- flow-through select operator MUX_3909_inst
    IMB39_3910 <= IMA79_3110 when (BITSEL_u8_u1_3906_wire(0) /=  '0') else IMA78_3100;
    -- logger for split-operator MUX_3917_inst flow-through 
    process(IMB40_3918) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3917_inst:flowthrough inputs: " & " BITSEL_u8_u1_3914_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3914_wire) & " IMA81_3130 = "& Convert_SLV_To_Hex_String(IMA81_3130) & " IMA80_3120 = "& Convert_SLV_To_Hex_String(IMA80_3120) & " outputs:" & " IMB40_3918= "  & Convert_SLV_To_Hex_String(IMB40_3918));
      --
    end process; 
    -- flow-through select operator MUX_3917_inst
    IMB40_3918 <= IMA81_3130 when (BITSEL_u8_u1_3914_wire(0) /=  '0') else IMA80_3120;
    -- logger for split-operator MUX_3925_inst flow-through 
    process(IMB41_3926) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3925_inst:flowthrough inputs: " & " BITSEL_u8_u1_3922_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3922_wire) & " IMA83_3150 = "& Convert_SLV_To_Hex_String(IMA83_3150) & " IMA82_3140 = "& Convert_SLV_To_Hex_String(IMA82_3140) & " outputs:" & " IMB41_3926= "  & Convert_SLV_To_Hex_String(IMB41_3926));
      --
    end process; 
    -- flow-through select operator MUX_3925_inst
    IMB41_3926 <= IMA83_3150 when (BITSEL_u8_u1_3922_wire(0) /=  '0') else IMA82_3140;
    -- logger for split-operator MUX_3933_inst flow-through 
    process(IMB42_3934) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3933_inst:flowthrough inputs: " & " BITSEL_u8_u1_3930_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3930_wire) & " IMA85_3170 = "& Convert_SLV_To_Hex_String(IMA85_3170) & " IMA84_3160 = "& Convert_SLV_To_Hex_String(IMA84_3160) & " outputs:" & " IMB42_3934= "  & Convert_SLV_To_Hex_String(IMB42_3934));
      --
    end process; 
    -- flow-through select operator MUX_3933_inst
    IMB42_3934 <= IMA85_3170 when (BITSEL_u8_u1_3930_wire(0) /=  '0') else IMA84_3160;
    -- logger for split-operator MUX_3941_inst flow-through 
    process(IMB43_3942) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3941_inst:flowthrough inputs: " & " BITSEL_u8_u1_3938_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3938_wire) & " IMA87_3190 = "& Convert_SLV_To_Hex_String(IMA87_3190) & " IMA86_3180 = "& Convert_SLV_To_Hex_String(IMA86_3180) & " outputs:" & " IMB43_3942= "  & Convert_SLV_To_Hex_String(IMB43_3942));
      --
    end process; 
    -- flow-through select operator MUX_3941_inst
    IMB43_3942 <= IMA87_3190 when (BITSEL_u8_u1_3938_wire(0) /=  '0') else IMA86_3180;
    -- logger for split-operator MUX_3949_inst flow-through 
    process(IMB44_3950) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3949_inst:flowthrough inputs: " & " BITSEL_u8_u1_3946_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3946_wire) & " IMA89_3210 = "& Convert_SLV_To_Hex_String(IMA89_3210) & " IMA88_3200 = "& Convert_SLV_To_Hex_String(IMA88_3200) & " outputs:" & " IMB44_3950= "  & Convert_SLV_To_Hex_String(IMB44_3950));
      --
    end process; 
    -- flow-through select operator MUX_3949_inst
    IMB44_3950 <= IMA89_3210 when (BITSEL_u8_u1_3946_wire(0) /=  '0') else IMA88_3200;
    -- logger for split-operator MUX_3957_inst flow-through 
    process(IMB45_3958) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3957_inst:flowthrough inputs: " & " BITSEL_u8_u1_3954_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3954_wire) & " IMA91_3230 = "& Convert_SLV_To_Hex_String(IMA91_3230) & " IMA90_3220 = "& Convert_SLV_To_Hex_String(IMA90_3220) & " outputs:" & " IMB45_3958= "  & Convert_SLV_To_Hex_String(IMB45_3958));
      --
    end process; 
    -- flow-through select operator MUX_3957_inst
    IMB45_3958 <= IMA91_3230 when (BITSEL_u8_u1_3954_wire(0) /=  '0') else IMA90_3220;
    -- logger for split-operator MUX_3965_inst flow-through 
    process(IMB46_3966) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3965_inst:flowthrough inputs: " & " BITSEL_u8_u1_3962_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3962_wire) & " IMA93_3250 = "& Convert_SLV_To_Hex_String(IMA93_3250) & " IMA92_3240 = "& Convert_SLV_To_Hex_String(IMA92_3240) & " outputs:" & " IMB46_3966= "  & Convert_SLV_To_Hex_String(IMB46_3966));
      --
    end process; 
    -- flow-through select operator MUX_3965_inst
    IMB46_3966 <= IMA93_3250 when (BITSEL_u8_u1_3962_wire(0) /=  '0') else IMA92_3240;
    -- logger for split-operator MUX_3973_inst flow-through 
    process(IMB47_3974) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3973_inst:flowthrough inputs: " & " BITSEL_u8_u1_3970_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3970_wire) & " IMA95_3270 = "& Convert_SLV_To_Hex_String(IMA95_3270) & " IMA94_3260 = "& Convert_SLV_To_Hex_String(IMA94_3260) & " outputs:" & " IMB47_3974= "  & Convert_SLV_To_Hex_String(IMB47_3974));
      --
    end process; 
    -- flow-through select operator MUX_3973_inst
    IMB47_3974 <= IMA95_3270 when (BITSEL_u8_u1_3970_wire(0) /=  '0') else IMA94_3260;
    -- logger for split-operator MUX_3981_inst flow-through 
    process(IMB48_3982) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3981_inst:flowthrough inputs: " & " BITSEL_u8_u1_3978_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3978_wire) & " IMA97_3290 = "& Convert_SLV_To_Hex_String(IMA97_3290) & " IMA96_3280 = "& Convert_SLV_To_Hex_String(IMA96_3280) & " outputs:" & " IMB48_3982= "  & Convert_SLV_To_Hex_String(IMB48_3982));
      --
    end process; 
    -- flow-through select operator MUX_3981_inst
    IMB48_3982 <= IMA97_3290 when (BITSEL_u8_u1_3978_wire(0) /=  '0') else IMA96_3280;
    -- logger for split-operator MUX_3989_inst flow-through 
    process(IMB49_3990) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3989_inst:flowthrough inputs: " & " BITSEL_u8_u1_3986_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3986_wire) & " IMA99_3310 = "& Convert_SLV_To_Hex_String(IMA99_3310) & " IMA98_3300 = "& Convert_SLV_To_Hex_String(IMA98_3300) & " outputs:" & " IMB49_3990= "  & Convert_SLV_To_Hex_String(IMB49_3990));
      --
    end process; 
    -- flow-through select operator MUX_3989_inst
    IMB49_3990 <= IMA99_3310 when (BITSEL_u8_u1_3986_wire(0) /=  '0') else IMA98_3300;
    -- logger for split-operator MUX_3997_inst flow-through 
    process(IMB50_3998) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_3997_inst:flowthrough inputs: " & " BITSEL_u8_u1_3994_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_3994_wire) & " IMA101_3330 = "& Convert_SLV_To_Hex_String(IMA101_3330) & " IMA100_3320 = "& Convert_SLV_To_Hex_String(IMA100_3320) & " outputs:" & " IMB50_3998= "  & Convert_SLV_To_Hex_String(IMB50_3998));
      --
    end process; 
    -- flow-through select operator MUX_3997_inst
    IMB50_3998 <= IMA101_3330 when (BITSEL_u8_u1_3994_wire(0) /=  '0') else IMA100_3320;
    -- logger for split-operator MUX_4005_inst flow-through 
    process(IMB51_4006) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_4005_inst:flowthrough inputs: " & " BITSEL_u8_u1_4002_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4002_wire) & " IMA103_3350 = "& Convert_SLV_To_Hex_String(IMA103_3350) & " IMA102_3340 = "& Convert_SLV_To_Hex_String(IMA102_3340) & " outputs:" & " IMB51_4006= "  & Convert_SLV_To_Hex_String(IMB51_4006));
      --
    end process; 
    -- flow-through select operator MUX_4005_inst
    IMB51_4006 <= IMA103_3350 when (BITSEL_u8_u1_4002_wire(0) /=  '0') else IMA102_3340;
    -- logger for split-operator MUX_4013_inst flow-through 
    process(IMB52_4014) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_4013_inst:flowthrough inputs: " & " BITSEL_u8_u1_4010_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4010_wire) & " IMA105_3370 = "& Convert_SLV_To_Hex_String(IMA105_3370) & " IMA104_3360 = "& Convert_SLV_To_Hex_String(IMA104_3360) & " outputs:" & " IMB52_4014= "  & Convert_SLV_To_Hex_String(IMB52_4014));
      --
    end process; 
    -- flow-through select operator MUX_4013_inst
    IMB52_4014 <= IMA105_3370 when (BITSEL_u8_u1_4010_wire(0) /=  '0') else IMA104_3360;
    -- logger for split-operator MUX_4021_inst flow-through 
    process(IMB53_4022) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_4021_inst:flowthrough inputs: " & " BITSEL_u8_u1_4018_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4018_wire) & " IMA107_3390 = "& Convert_SLV_To_Hex_String(IMA107_3390) & " IMA106_3380 = "& Convert_SLV_To_Hex_String(IMA106_3380) & " outputs:" & " IMB53_4022= "  & Convert_SLV_To_Hex_String(IMB53_4022));
      --
    end process; 
    -- flow-through select operator MUX_4021_inst
    IMB53_4022 <= IMA107_3390 when (BITSEL_u8_u1_4018_wire(0) /=  '0') else IMA106_3380;
    -- logger for split-operator MUX_4029_inst flow-through 
    process(IMB54_4030) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_4029_inst:flowthrough inputs: " & " BITSEL_u8_u1_4026_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4026_wire) & " IMA109_3410 = "& Convert_SLV_To_Hex_String(IMA109_3410) & " IMA108_3400 = "& Convert_SLV_To_Hex_String(IMA108_3400) & " outputs:" & " IMB54_4030= "  & Convert_SLV_To_Hex_String(IMB54_4030));
      --
    end process; 
    -- flow-through select operator MUX_4029_inst
    IMB54_4030 <= IMA109_3410 when (BITSEL_u8_u1_4026_wire(0) /=  '0') else IMA108_3400;
    -- logger for split-operator MUX_4037_inst flow-through 
    process(IMB55_4038) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_4037_inst:flowthrough inputs: " & " BITSEL_u8_u1_4034_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4034_wire) & " IMA111_3430 = "& Convert_SLV_To_Hex_String(IMA111_3430) & " IMA110_3420 = "& Convert_SLV_To_Hex_String(IMA110_3420) & " outputs:" & " IMB55_4038= "  & Convert_SLV_To_Hex_String(IMB55_4038));
      --
    end process; 
    -- flow-through select operator MUX_4037_inst
    IMB55_4038 <= IMA111_3430 when (BITSEL_u8_u1_4034_wire(0) /=  '0') else IMA110_3420;
    -- logger for split-operator MUX_4045_inst flow-through 
    process(IMB56_4046) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_4045_inst:flowthrough inputs: " & " BITSEL_u8_u1_4042_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4042_wire) & " IMA113_3450 = "& Convert_SLV_To_Hex_String(IMA113_3450) & " IMA112_3440 = "& Convert_SLV_To_Hex_String(IMA112_3440) & " outputs:" & " IMB56_4046= "  & Convert_SLV_To_Hex_String(IMB56_4046));
      --
    end process; 
    -- flow-through select operator MUX_4045_inst
    IMB56_4046 <= IMA113_3450 when (BITSEL_u8_u1_4042_wire(0) /=  '0') else IMA112_3440;
    -- logger for split-operator MUX_4053_inst flow-through 
    process(IMB57_4054) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_4053_inst:flowthrough inputs: " & " BITSEL_u8_u1_4050_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4050_wire) & " IMA115_3470 = "& Convert_SLV_To_Hex_String(IMA115_3470) & " IMA114_3460 = "& Convert_SLV_To_Hex_String(IMA114_3460) & " outputs:" & " IMB57_4054= "  & Convert_SLV_To_Hex_String(IMB57_4054));
      --
    end process; 
    -- flow-through select operator MUX_4053_inst
    IMB57_4054 <= IMA115_3470 when (BITSEL_u8_u1_4050_wire(0) /=  '0') else IMA114_3460;
    -- logger for split-operator MUX_4061_inst flow-through 
    process(IMB58_4062) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_4061_inst:flowthrough inputs: " & " BITSEL_u8_u1_4058_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4058_wire) & " IMA117_3490 = "& Convert_SLV_To_Hex_String(IMA117_3490) & " IMA116_3480 = "& Convert_SLV_To_Hex_String(IMA116_3480) & " outputs:" & " IMB58_4062= "  & Convert_SLV_To_Hex_String(IMB58_4062));
      --
    end process; 
    -- flow-through select operator MUX_4061_inst
    IMB58_4062 <= IMA117_3490 when (BITSEL_u8_u1_4058_wire(0) /=  '0') else IMA116_3480;
    -- logger for split-operator MUX_4069_inst flow-through 
    process(IMB59_4070) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_4069_inst:flowthrough inputs: " & " BITSEL_u8_u1_4066_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4066_wire) & " IMA119_3510 = "& Convert_SLV_To_Hex_String(IMA119_3510) & " IMA118_3500 = "& Convert_SLV_To_Hex_String(IMA118_3500) & " outputs:" & " IMB59_4070= "  & Convert_SLV_To_Hex_String(IMB59_4070));
      --
    end process; 
    -- flow-through select operator MUX_4069_inst
    IMB59_4070 <= IMA119_3510 when (BITSEL_u8_u1_4066_wire(0) /=  '0') else IMA118_3500;
    -- logger for split-operator MUX_4077_inst flow-through 
    process(IMB60_4078) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_4077_inst:flowthrough inputs: " & " BITSEL_u8_u1_4074_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4074_wire) & " IMA121_3530 = "& Convert_SLV_To_Hex_String(IMA121_3530) & " IMA120_3520 = "& Convert_SLV_To_Hex_String(IMA120_3520) & " outputs:" & " IMB60_4078= "  & Convert_SLV_To_Hex_String(IMB60_4078));
      --
    end process; 
    -- flow-through select operator MUX_4077_inst
    IMB60_4078 <= IMA121_3530 when (BITSEL_u8_u1_4074_wire(0) /=  '0') else IMA120_3520;
    -- logger for split-operator MUX_4085_inst flow-through 
    process(IMB61_4086) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_4085_inst:flowthrough inputs: " & " BITSEL_u8_u1_4082_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4082_wire) & " IMA123_3550 = "& Convert_SLV_To_Hex_String(IMA123_3550) & " IMA122_3540 = "& Convert_SLV_To_Hex_String(IMA122_3540) & " outputs:" & " IMB61_4086= "  & Convert_SLV_To_Hex_String(IMB61_4086));
      --
    end process; 
    -- flow-through select operator MUX_4085_inst
    IMB61_4086 <= IMA123_3550 when (BITSEL_u8_u1_4082_wire(0) /=  '0') else IMA122_3540;
    -- logger for split-operator MUX_4093_inst flow-through 
    process(IMB62_4094) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_4093_inst:flowthrough inputs: " & " BITSEL_u8_u1_4090_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4090_wire) & " IMA125_3570 = "& Convert_SLV_To_Hex_String(IMA125_3570) & " IMA124_3560 = "& Convert_SLV_To_Hex_String(IMA124_3560) & " outputs:" & " IMB62_4094= "  & Convert_SLV_To_Hex_String(IMB62_4094));
      --
    end process; 
    -- flow-through select operator MUX_4093_inst
    IMB62_4094 <= IMA125_3570 when (BITSEL_u8_u1_4090_wire(0) /=  '0') else IMA124_3560;
    -- logger for split-operator MUX_4101_inst flow-through 
    process(IMB63_4102) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_4101_inst:flowthrough inputs: " & " BITSEL_u8_u1_4098_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4098_wire) & " IMA127_3590 = "& Convert_SLV_To_Hex_String(IMA127_3590) & " IMA126_3580 = "& Convert_SLV_To_Hex_String(IMA126_3580) & " outputs:" & " IMB63_4102= "  & Convert_SLV_To_Hex_String(IMB63_4102));
      --
    end process; 
    -- flow-through select operator MUX_4101_inst
    IMB63_4102 <= IMA127_3590 when (BITSEL_u8_u1_4098_wire(0) /=  '0') else IMA126_3580;
    -- logger for split-operator MUX_4109_inst flow-through 
    process(IMC0_4110) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_4109_inst:flowthrough inputs: " & " BITSEL_u8_u1_4106_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4106_wire) & " IMB1_3606 = "& Convert_SLV_To_Hex_String(IMB1_3606) & " IMB0_3598 = "& Convert_SLV_To_Hex_String(IMB0_3598) & " outputs:" & " IMC0_4110= "  & Convert_SLV_To_Hex_String(IMC0_4110));
      --
    end process; 
    -- flow-through select operator MUX_4109_inst
    IMC0_4110 <= IMB1_3606 when (BITSEL_u8_u1_4106_wire(0) /=  '0') else IMB0_3598;
    -- logger for split-operator MUX_4117_inst flow-through 
    process(IMC1_4118) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_4117_inst:flowthrough inputs: " & " BITSEL_u8_u1_4114_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4114_wire) & " IMB3_3622 = "& Convert_SLV_To_Hex_String(IMB3_3622) & " IMB2_3614 = "& Convert_SLV_To_Hex_String(IMB2_3614) & " outputs:" & " IMC1_4118= "  & Convert_SLV_To_Hex_String(IMC1_4118));
      --
    end process; 
    -- flow-through select operator MUX_4117_inst
    IMC1_4118 <= IMB3_3622 when (BITSEL_u8_u1_4114_wire(0) /=  '0') else IMB2_3614;
    -- logger for split-operator MUX_4125_inst flow-through 
    process(IMC2_4126) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_4125_inst:flowthrough inputs: " & " BITSEL_u8_u1_4122_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4122_wire) & " IMB5_3638 = "& Convert_SLV_To_Hex_String(IMB5_3638) & " IMB4_3630 = "& Convert_SLV_To_Hex_String(IMB4_3630) & " outputs:" & " IMC2_4126= "  & Convert_SLV_To_Hex_String(IMC2_4126));
      --
    end process; 
    -- flow-through select operator MUX_4125_inst
    IMC2_4126 <= IMB5_3638 when (BITSEL_u8_u1_4122_wire(0) /=  '0') else IMB4_3630;
    -- logger for split-operator MUX_4133_inst flow-through 
    process(IMC3_4134) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_4133_inst:flowthrough inputs: " & " BITSEL_u8_u1_4130_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4130_wire) & " IMB7_3654 = "& Convert_SLV_To_Hex_String(IMB7_3654) & " IMB6_3646 = "& Convert_SLV_To_Hex_String(IMB6_3646) & " outputs:" & " IMC3_4134= "  & Convert_SLV_To_Hex_String(IMC3_4134));
      --
    end process; 
    -- flow-through select operator MUX_4133_inst
    IMC3_4134 <= IMB7_3654 when (BITSEL_u8_u1_4130_wire(0) /=  '0') else IMB6_3646;
    -- logger for split-operator MUX_4141_inst flow-through 
    process(IMC4_4142) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_4141_inst:flowthrough inputs: " & " BITSEL_u8_u1_4138_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4138_wire) & " IMB9_3670 = "& Convert_SLV_To_Hex_String(IMB9_3670) & " IMB8_3662 = "& Convert_SLV_To_Hex_String(IMB8_3662) & " outputs:" & " IMC4_4142= "  & Convert_SLV_To_Hex_String(IMC4_4142));
      --
    end process; 
    -- flow-through select operator MUX_4141_inst
    IMC4_4142 <= IMB9_3670 when (BITSEL_u8_u1_4138_wire(0) /=  '0') else IMB8_3662;
    -- logger for split-operator MUX_4149_inst flow-through 
    process(IMC5_4150) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_4149_inst:flowthrough inputs: " & " BITSEL_u8_u1_4146_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4146_wire) & " IMB11_3686 = "& Convert_SLV_To_Hex_String(IMB11_3686) & " IMB10_3678 = "& Convert_SLV_To_Hex_String(IMB10_3678) & " outputs:" & " IMC5_4150= "  & Convert_SLV_To_Hex_String(IMC5_4150));
      --
    end process; 
    -- flow-through select operator MUX_4149_inst
    IMC5_4150 <= IMB11_3686 when (BITSEL_u8_u1_4146_wire(0) /=  '0') else IMB10_3678;
    -- logger for split-operator MUX_4157_inst flow-through 
    process(IMC6_4158) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_4157_inst:flowthrough inputs: " & " BITSEL_u8_u1_4154_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4154_wire) & " IMB13_3702 = "& Convert_SLV_To_Hex_String(IMB13_3702) & " IMB12_3694 = "& Convert_SLV_To_Hex_String(IMB12_3694) & " outputs:" & " IMC6_4158= "  & Convert_SLV_To_Hex_String(IMC6_4158));
      --
    end process; 
    -- flow-through select operator MUX_4157_inst
    IMC6_4158 <= IMB13_3702 when (BITSEL_u8_u1_4154_wire(0) /=  '0') else IMB12_3694;
    -- logger for split-operator MUX_4165_inst flow-through 
    process(IMC7_4166) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_4165_inst:flowthrough inputs: " & " BITSEL_u8_u1_4162_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4162_wire) & " IMB15_3718 = "& Convert_SLV_To_Hex_String(IMB15_3718) & " IMB14_3710 = "& Convert_SLV_To_Hex_String(IMB14_3710) & " outputs:" & " IMC7_4166= "  & Convert_SLV_To_Hex_String(IMC7_4166));
      --
    end process; 
    -- flow-through select operator MUX_4165_inst
    IMC7_4166 <= IMB15_3718 when (BITSEL_u8_u1_4162_wire(0) /=  '0') else IMB14_3710;
    -- logger for split-operator MUX_4173_inst flow-through 
    process(IMC8_4174) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_4173_inst:flowthrough inputs: " & " BITSEL_u8_u1_4170_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4170_wire) & " IMB17_3734 = "& Convert_SLV_To_Hex_String(IMB17_3734) & " IMB16_3726 = "& Convert_SLV_To_Hex_String(IMB16_3726) & " outputs:" & " IMC8_4174= "  & Convert_SLV_To_Hex_String(IMC8_4174));
      --
    end process; 
    -- flow-through select operator MUX_4173_inst
    IMC8_4174 <= IMB17_3734 when (BITSEL_u8_u1_4170_wire(0) /=  '0') else IMB16_3726;
    -- logger for split-operator MUX_4181_inst flow-through 
    process(IMC9_4182) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_4181_inst:flowthrough inputs: " & " BITSEL_u8_u1_4178_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4178_wire) & " IMB19_3750 = "& Convert_SLV_To_Hex_String(IMB19_3750) & " IMB18_3742 = "& Convert_SLV_To_Hex_String(IMB18_3742) & " outputs:" & " IMC9_4182= "  & Convert_SLV_To_Hex_String(IMC9_4182));
      --
    end process; 
    -- flow-through select operator MUX_4181_inst
    IMC9_4182 <= IMB19_3750 when (BITSEL_u8_u1_4178_wire(0) /=  '0') else IMB18_3742;
    -- logger for split-operator MUX_4189_inst flow-through 
    process(IMC10_4190) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_4189_inst:flowthrough inputs: " & " BITSEL_u8_u1_4186_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4186_wire) & " IMB21_3766 = "& Convert_SLV_To_Hex_String(IMB21_3766) & " IMB20_3758 = "& Convert_SLV_To_Hex_String(IMB20_3758) & " outputs:" & " IMC10_4190= "  & Convert_SLV_To_Hex_String(IMC10_4190));
      --
    end process; 
    -- flow-through select operator MUX_4189_inst
    IMC10_4190 <= IMB21_3766 when (BITSEL_u8_u1_4186_wire(0) /=  '0') else IMB20_3758;
    -- logger for split-operator MUX_4197_inst flow-through 
    process(IMC11_4198) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_4197_inst:flowthrough inputs: " & " BITSEL_u8_u1_4194_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4194_wire) & " IMB23_3782 = "& Convert_SLV_To_Hex_String(IMB23_3782) & " IMB22_3774 = "& Convert_SLV_To_Hex_String(IMB22_3774) & " outputs:" & " IMC11_4198= "  & Convert_SLV_To_Hex_String(IMC11_4198));
      --
    end process; 
    -- flow-through select operator MUX_4197_inst
    IMC11_4198 <= IMB23_3782 when (BITSEL_u8_u1_4194_wire(0) /=  '0') else IMB22_3774;
    -- logger for split-operator MUX_4205_inst flow-through 
    process(IMC12_4206) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_4205_inst:flowthrough inputs: " & " BITSEL_u8_u1_4202_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4202_wire) & " IMB25_3798 = "& Convert_SLV_To_Hex_String(IMB25_3798) & " IMB24_3790 = "& Convert_SLV_To_Hex_String(IMB24_3790) & " outputs:" & " IMC12_4206= "  & Convert_SLV_To_Hex_String(IMC12_4206));
      --
    end process; 
    -- flow-through select operator MUX_4205_inst
    IMC12_4206 <= IMB25_3798 when (BITSEL_u8_u1_4202_wire(0) /=  '0') else IMB24_3790;
    -- logger for split-operator MUX_4213_inst flow-through 
    process(IMC13_4214) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_4213_inst:flowthrough inputs: " & " BITSEL_u8_u1_4210_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4210_wire) & " IMB27_3814 = "& Convert_SLV_To_Hex_String(IMB27_3814) & " IMB26_3806 = "& Convert_SLV_To_Hex_String(IMB26_3806) & " outputs:" & " IMC13_4214= "  & Convert_SLV_To_Hex_String(IMC13_4214));
      --
    end process; 
    -- flow-through select operator MUX_4213_inst
    IMC13_4214 <= IMB27_3814 when (BITSEL_u8_u1_4210_wire(0) /=  '0') else IMB26_3806;
    -- logger for split-operator MUX_4221_inst flow-through 
    process(IMC14_4222) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_4221_inst:flowthrough inputs: " & " BITSEL_u8_u1_4218_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4218_wire) & " IMB29_3830 = "& Convert_SLV_To_Hex_String(IMB29_3830) & " IMB28_3822 = "& Convert_SLV_To_Hex_String(IMB28_3822) & " outputs:" & " IMC14_4222= "  & Convert_SLV_To_Hex_String(IMC14_4222));
      --
    end process; 
    -- flow-through select operator MUX_4221_inst
    IMC14_4222 <= IMB29_3830 when (BITSEL_u8_u1_4218_wire(0) /=  '0') else IMB28_3822;
    -- logger for split-operator MUX_4229_inst flow-through 
    process(IMC15_4230) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_4229_inst:flowthrough inputs: " & " BITSEL_u8_u1_4226_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4226_wire) & " IMB31_3846 = "& Convert_SLV_To_Hex_String(IMB31_3846) & " IMB30_3838 = "& Convert_SLV_To_Hex_String(IMB30_3838) & " outputs:" & " IMC15_4230= "  & Convert_SLV_To_Hex_String(IMC15_4230));
      --
    end process; 
    -- flow-through select operator MUX_4229_inst
    IMC15_4230 <= IMB31_3846 when (BITSEL_u8_u1_4226_wire(0) /=  '0') else IMB30_3838;
    -- logger for split-operator MUX_4237_inst flow-through 
    process(IMC16_4238) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_4237_inst:flowthrough inputs: " & " BITSEL_u8_u1_4234_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4234_wire) & " IMB33_3862 = "& Convert_SLV_To_Hex_String(IMB33_3862) & " IMB32_3854 = "& Convert_SLV_To_Hex_String(IMB32_3854) & " outputs:" & " IMC16_4238= "  & Convert_SLV_To_Hex_String(IMC16_4238));
      --
    end process; 
    -- flow-through select operator MUX_4237_inst
    IMC16_4238 <= IMB33_3862 when (BITSEL_u8_u1_4234_wire(0) /=  '0') else IMB32_3854;
    -- logger for split-operator MUX_4245_inst flow-through 
    process(IMC17_4246) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_4245_inst:flowthrough inputs: " & " BITSEL_u8_u1_4242_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4242_wire) & " IMB35_3878 = "& Convert_SLV_To_Hex_String(IMB35_3878) & " IMB34_3870 = "& Convert_SLV_To_Hex_String(IMB34_3870) & " outputs:" & " IMC17_4246= "  & Convert_SLV_To_Hex_String(IMC17_4246));
      --
    end process; 
    -- flow-through select operator MUX_4245_inst
    IMC17_4246 <= IMB35_3878 when (BITSEL_u8_u1_4242_wire(0) /=  '0') else IMB34_3870;
    -- logger for split-operator MUX_4253_inst flow-through 
    process(IMC18_4254) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_4253_inst:flowthrough inputs: " & " BITSEL_u8_u1_4250_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4250_wire) & " IMB37_3894 = "& Convert_SLV_To_Hex_String(IMB37_3894) & " IMB36_3886 = "& Convert_SLV_To_Hex_String(IMB36_3886) & " outputs:" & " IMC18_4254= "  & Convert_SLV_To_Hex_String(IMC18_4254));
      --
    end process; 
    -- flow-through select operator MUX_4253_inst
    IMC18_4254 <= IMB37_3894 when (BITSEL_u8_u1_4250_wire(0) /=  '0') else IMB36_3886;
    -- logger for split-operator MUX_4261_inst flow-through 
    process(IMC19_4262) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_4261_inst:flowthrough inputs: " & " BITSEL_u8_u1_4258_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4258_wire) & " IMB39_3910 = "& Convert_SLV_To_Hex_String(IMB39_3910) & " IMB38_3902 = "& Convert_SLV_To_Hex_String(IMB38_3902) & " outputs:" & " IMC19_4262= "  & Convert_SLV_To_Hex_String(IMC19_4262));
      --
    end process; 
    -- flow-through select operator MUX_4261_inst
    IMC19_4262 <= IMB39_3910 when (BITSEL_u8_u1_4258_wire(0) /=  '0') else IMB38_3902;
    -- logger for split-operator MUX_4269_inst flow-through 
    process(IMC20_4270) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_4269_inst:flowthrough inputs: " & " BITSEL_u8_u1_4266_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4266_wire) & " IMB41_3926 = "& Convert_SLV_To_Hex_String(IMB41_3926) & " IMB40_3918 = "& Convert_SLV_To_Hex_String(IMB40_3918) & " outputs:" & " IMC20_4270= "  & Convert_SLV_To_Hex_String(IMC20_4270));
      --
    end process; 
    -- flow-through select operator MUX_4269_inst
    IMC20_4270 <= IMB41_3926 when (BITSEL_u8_u1_4266_wire(0) /=  '0') else IMB40_3918;
    -- logger for split-operator MUX_4277_inst flow-through 
    process(IMC21_4278) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_4277_inst:flowthrough inputs: " & " BITSEL_u8_u1_4274_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4274_wire) & " IMB43_3942 = "& Convert_SLV_To_Hex_String(IMB43_3942) & " IMB42_3934 = "& Convert_SLV_To_Hex_String(IMB42_3934) & " outputs:" & " IMC21_4278= "  & Convert_SLV_To_Hex_String(IMC21_4278));
      --
    end process; 
    -- flow-through select operator MUX_4277_inst
    IMC21_4278 <= IMB43_3942 when (BITSEL_u8_u1_4274_wire(0) /=  '0') else IMB42_3934;
    -- logger for split-operator MUX_4285_inst flow-through 
    process(IMC22_4286) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_4285_inst:flowthrough inputs: " & " BITSEL_u8_u1_4282_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4282_wire) & " IMB45_3958 = "& Convert_SLV_To_Hex_String(IMB45_3958) & " IMB44_3950 = "& Convert_SLV_To_Hex_String(IMB44_3950) & " outputs:" & " IMC22_4286= "  & Convert_SLV_To_Hex_String(IMC22_4286));
      --
    end process; 
    -- flow-through select operator MUX_4285_inst
    IMC22_4286 <= IMB45_3958 when (BITSEL_u8_u1_4282_wire(0) /=  '0') else IMB44_3950;
    -- logger for split-operator MUX_4293_inst flow-through 
    process(IMC23_4294) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_4293_inst:flowthrough inputs: " & " BITSEL_u8_u1_4290_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4290_wire) & " IMB47_3974 = "& Convert_SLV_To_Hex_String(IMB47_3974) & " IMB46_3966 = "& Convert_SLV_To_Hex_String(IMB46_3966) & " outputs:" & " IMC23_4294= "  & Convert_SLV_To_Hex_String(IMC23_4294));
      --
    end process; 
    -- flow-through select operator MUX_4293_inst
    IMC23_4294 <= IMB47_3974 when (BITSEL_u8_u1_4290_wire(0) /=  '0') else IMB46_3966;
    -- logger for split-operator MUX_4301_inst flow-through 
    process(IMC24_4302) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_4301_inst:flowthrough inputs: " & " BITSEL_u8_u1_4298_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4298_wire) & " IMB49_3990 = "& Convert_SLV_To_Hex_String(IMB49_3990) & " IMB48_3982 = "& Convert_SLV_To_Hex_String(IMB48_3982) & " outputs:" & " IMC24_4302= "  & Convert_SLV_To_Hex_String(IMC24_4302));
      --
    end process; 
    -- flow-through select operator MUX_4301_inst
    IMC24_4302 <= IMB49_3990 when (BITSEL_u8_u1_4298_wire(0) /=  '0') else IMB48_3982;
    -- logger for split-operator MUX_4309_inst flow-through 
    process(IMC25_4310) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_4309_inst:flowthrough inputs: " & " BITSEL_u8_u1_4306_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4306_wire) & " IMB51_4006 = "& Convert_SLV_To_Hex_String(IMB51_4006) & " IMB50_3998 = "& Convert_SLV_To_Hex_String(IMB50_3998) & " outputs:" & " IMC25_4310= "  & Convert_SLV_To_Hex_String(IMC25_4310));
      --
    end process; 
    -- flow-through select operator MUX_4309_inst
    IMC25_4310 <= IMB51_4006 when (BITSEL_u8_u1_4306_wire(0) /=  '0') else IMB50_3998;
    -- logger for split-operator MUX_4317_inst flow-through 
    process(IMC26_4318) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_4317_inst:flowthrough inputs: " & " BITSEL_u8_u1_4314_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4314_wire) & " IMB53_4022 = "& Convert_SLV_To_Hex_String(IMB53_4022) & " IMB52_4014 = "& Convert_SLV_To_Hex_String(IMB52_4014) & " outputs:" & " IMC26_4318= "  & Convert_SLV_To_Hex_String(IMC26_4318));
      --
    end process; 
    -- flow-through select operator MUX_4317_inst
    IMC26_4318 <= IMB53_4022 when (BITSEL_u8_u1_4314_wire(0) /=  '0') else IMB52_4014;
    -- logger for split-operator MUX_4325_inst flow-through 
    process(IMC27_4326) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_4325_inst:flowthrough inputs: " & " BITSEL_u8_u1_4322_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4322_wire) & " IMB55_4038 = "& Convert_SLV_To_Hex_String(IMB55_4038) & " IMB54_4030 = "& Convert_SLV_To_Hex_String(IMB54_4030) & " outputs:" & " IMC27_4326= "  & Convert_SLV_To_Hex_String(IMC27_4326));
      --
    end process; 
    -- flow-through select operator MUX_4325_inst
    IMC27_4326 <= IMB55_4038 when (BITSEL_u8_u1_4322_wire(0) /=  '0') else IMB54_4030;
    -- logger for split-operator MUX_4333_inst flow-through 
    process(IMC28_4334) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_4333_inst:flowthrough inputs: " & " BITSEL_u8_u1_4330_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4330_wire) & " IMB57_4054 = "& Convert_SLV_To_Hex_String(IMB57_4054) & " IMB56_4046 = "& Convert_SLV_To_Hex_String(IMB56_4046) & " outputs:" & " IMC28_4334= "  & Convert_SLV_To_Hex_String(IMC28_4334));
      --
    end process; 
    -- flow-through select operator MUX_4333_inst
    IMC28_4334 <= IMB57_4054 when (BITSEL_u8_u1_4330_wire(0) /=  '0') else IMB56_4046;
    -- logger for split-operator MUX_4341_inst flow-through 
    process(IMC29_4342) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_4341_inst:flowthrough inputs: " & " BITSEL_u8_u1_4338_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4338_wire) & " IMB59_4070 = "& Convert_SLV_To_Hex_String(IMB59_4070) & " IMB58_4062 = "& Convert_SLV_To_Hex_String(IMB58_4062) & " outputs:" & " IMC29_4342= "  & Convert_SLV_To_Hex_String(IMC29_4342));
      --
    end process; 
    -- flow-through select operator MUX_4341_inst
    IMC29_4342 <= IMB59_4070 when (BITSEL_u8_u1_4338_wire(0) /=  '0') else IMB58_4062;
    -- logger for split-operator MUX_4349_inst flow-through 
    process(IMC30_4350) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_4349_inst:flowthrough inputs: " & " BITSEL_u8_u1_4346_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4346_wire) & " IMB61_4086 = "& Convert_SLV_To_Hex_String(IMB61_4086) & " IMB60_4078 = "& Convert_SLV_To_Hex_String(IMB60_4078) & " outputs:" & " IMC30_4350= "  & Convert_SLV_To_Hex_String(IMC30_4350));
      --
    end process; 
    -- flow-through select operator MUX_4349_inst
    IMC30_4350 <= IMB61_4086 when (BITSEL_u8_u1_4346_wire(0) /=  '0') else IMB60_4078;
    -- logger for split-operator MUX_4357_inst flow-through 
    process(IMC31_4358) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_4357_inst:flowthrough inputs: " & " BITSEL_u8_u1_4354_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4354_wire) & " IMB63_4102 = "& Convert_SLV_To_Hex_String(IMB63_4102) & " IMB62_4094 = "& Convert_SLV_To_Hex_String(IMB62_4094) & " outputs:" & " IMC31_4358= "  & Convert_SLV_To_Hex_String(IMC31_4358));
      --
    end process; 
    -- flow-through select operator MUX_4357_inst
    IMC31_4358 <= IMB63_4102 when (BITSEL_u8_u1_4354_wire(0) /=  '0') else IMB62_4094;
    -- logger for split-operator MUX_4365_inst flow-through 
    process(IMD0_4366) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_4365_inst:flowthrough inputs: " & " BITSEL_u8_u1_4362_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4362_wire) & " IMC1_4118 = "& Convert_SLV_To_Hex_String(IMC1_4118) & " IMC0_4110 = "& Convert_SLV_To_Hex_String(IMC0_4110) & " outputs:" & " IMD0_4366= "  & Convert_SLV_To_Hex_String(IMD0_4366));
      --
    end process; 
    -- flow-through select operator MUX_4365_inst
    IMD0_4366 <= IMC1_4118 when (BITSEL_u8_u1_4362_wire(0) /=  '0') else IMC0_4110;
    -- logger for split-operator MUX_4373_inst flow-through 
    process(IMD1_4374) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_4373_inst:flowthrough inputs: " & " BITSEL_u8_u1_4370_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4370_wire) & " IMC3_4134 = "& Convert_SLV_To_Hex_String(IMC3_4134) & " IMC2_4126 = "& Convert_SLV_To_Hex_String(IMC2_4126) & " outputs:" & " IMD1_4374= "  & Convert_SLV_To_Hex_String(IMD1_4374));
      --
    end process; 
    -- flow-through select operator MUX_4373_inst
    IMD1_4374 <= IMC3_4134 when (BITSEL_u8_u1_4370_wire(0) /=  '0') else IMC2_4126;
    -- logger for split-operator MUX_4381_inst flow-through 
    process(IMD2_4382) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_4381_inst:flowthrough inputs: " & " BITSEL_u8_u1_4378_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4378_wire) & " IMC5_4150 = "& Convert_SLV_To_Hex_String(IMC5_4150) & " IMC4_4142 = "& Convert_SLV_To_Hex_String(IMC4_4142) & " outputs:" & " IMD2_4382= "  & Convert_SLV_To_Hex_String(IMD2_4382));
      --
    end process; 
    -- flow-through select operator MUX_4381_inst
    IMD2_4382 <= IMC5_4150 when (BITSEL_u8_u1_4378_wire(0) /=  '0') else IMC4_4142;
    -- logger for split-operator MUX_4389_inst flow-through 
    process(IMD3_4390) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_4389_inst:flowthrough inputs: " & " BITSEL_u8_u1_4386_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4386_wire) & " IMC7_4166 = "& Convert_SLV_To_Hex_String(IMC7_4166) & " IMC6_4158 = "& Convert_SLV_To_Hex_String(IMC6_4158) & " outputs:" & " IMD3_4390= "  & Convert_SLV_To_Hex_String(IMD3_4390));
      --
    end process; 
    -- flow-through select operator MUX_4389_inst
    IMD3_4390 <= IMC7_4166 when (BITSEL_u8_u1_4386_wire(0) /=  '0') else IMC6_4158;
    -- logger for split-operator MUX_4397_inst flow-through 
    process(IMD4_4398) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_4397_inst:flowthrough inputs: " & " BITSEL_u8_u1_4394_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4394_wire) & " IMC9_4182 = "& Convert_SLV_To_Hex_String(IMC9_4182) & " IMC8_4174 = "& Convert_SLV_To_Hex_String(IMC8_4174) & " outputs:" & " IMD4_4398= "  & Convert_SLV_To_Hex_String(IMD4_4398));
      --
    end process; 
    -- flow-through select operator MUX_4397_inst
    IMD4_4398 <= IMC9_4182 when (BITSEL_u8_u1_4394_wire(0) /=  '0') else IMC8_4174;
    -- logger for split-operator MUX_4405_inst flow-through 
    process(IMD5_4406) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_4405_inst:flowthrough inputs: " & " BITSEL_u8_u1_4402_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4402_wire) & " IMC11_4198 = "& Convert_SLV_To_Hex_String(IMC11_4198) & " IMC10_4190 = "& Convert_SLV_To_Hex_String(IMC10_4190) & " outputs:" & " IMD5_4406= "  & Convert_SLV_To_Hex_String(IMD5_4406));
      --
    end process; 
    -- flow-through select operator MUX_4405_inst
    IMD5_4406 <= IMC11_4198 when (BITSEL_u8_u1_4402_wire(0) /=  '0') else IMC10_4190;
    -- logger for split-operator MUX_4413_inst flow-through 
    process(IMD6_4414) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_4413_inst:flowthrough inputs: " & " BITSEL_u8_u1_4410_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4410_wire) & " IMC13_4214 = "& Convert_SLV_To_Hex_String(IMC13_4214) & " IMC12_4206 = "& Convert_SLV_To_Hex_String(IMC12_4206) & " outputs:" & " IMD6_4414= "  & Convert_SLV_To_Hex_String(IMD6_4414));
      --
    end process; 
    -- flow-through select operator MUX_4413_inst
    IMD6_4414 <= IMC13_4214 when (BITSEL_u8_u1_4410_wire(0) /=  '0') else IMC12_4206;
    -- logger for split-operator MUX_4421_inst flow-through 
    process(IMD7_4422) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_4421_inst:flowthrough inputs: " & " BITSEL_u8_u1_4418_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4418_wire) & " IMC15_4230 = "& Convert_SLV_To_Hex_String(IMC15_4230) & " IMC14_4222 = "& Convert_SLV_To_Hex_String(IMC14_4222) & " outputs:" & " IMD7_4422= "  & Convert_SLV_To_Hex_String(IMD7_4422));
      --
    end process; 
    -- flow-through select operator MUX_4421_inst
    IMD7_4422 <= IMC15_4230 when (BITSEL_u8_u1_4418_wire(0) /=  '0') else IMC14_4222;
    -- logger for split-operator MUX_4429_inst flow-through 
    process(IMD8_4430) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_4429_inst:flowthrough inputs: " & " BITSEL_u8_u1_4426_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4426_wire) & " IMC17_4246 = "& Convert_SLV_To_Hex_String(IMC17_4246) & " IMC16_4238 = "& Convert_SLV_To_Hex_String(IMC16_4238) & " outputs:" & " IMD8_4430= "  & Convert_SLV_To_Hex_String(IMD8_4430));
      --
    end process; 
    -- flow-through select operator MUX_4429_inst
    IMD8_4430 <= IMC17_4246 when (BITSEL_u8_u1_4426_wire(0) /=  '0') else IMC16_4238;
    -- logger for split-operator MUX_4437_inst flow-through 
    process(IMD9_4438) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_4437_inst:flowthrough inputs: " & " BITSEL_u8_u1_4434_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4434_wire) & " IMC19_4262 = "& Convert_SLV_To_Hex_String(IMC19_4262) & " IMC18_4254 = "& Convert_SLV_To_Hex_String(IMC18_4254) & " outputs:" & " IMD9_4438= "  & Convert_SLV_To_Hex_String(IMD9_4438));
      --
    end process; 
    -- flow-through select operator MUX_4437_inst
    IMD9_4438 <= IMC19_4262 when (BITSEL_u8_u1_4434_wire(0) /=  '0') else IMC18_4254;
    -- logger for split-operator MUX_4445_inst flow-through 
    process(IMD10_4446) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_4445_inst:flowthrough inputs: " & " BITSEL_u8_u1_4442_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4442_wire) & " IMC21_4278 = "& Convert_SLV_To_Hex_String(IMC21_4278) & " IMC20_4270 = "& Convert_SLV_To_Hex_String(IMC20_4270) & " outputs:" & " IMD10_4446= "  & Convert_SLV_To_Hex_String(IMD10_4446));
      --
    end process; 
    -- flow-through select operator MUX_4445_inst
    IMD10_4446 <= IMC21_4278 when (BITSEL_u8_u1_4442_wire(0) /=  '0') else IMC20_4270;
    -- logger for split-operator MUX_4453_inst flow-through 
    process(IMD11_4454) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_4453_inst:flowthrough inputs: " & " BITSEL_u8_u1_4450_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4450_wire) & " IMC23_4294 = "& Convert_SLV_To_Hex_String(IMC23_4294) & " IMC22_4286 = "& Convert_SLV_To_Hex_String(IMC22_4286) & " outputs:" & " IMD11_4454= "  & Convert_SLV_To_Hex_String(IMD11_4454));
      --
    end process; 
    -- flow-through select operator MUX_4453_inst
    IMD11_4454 <= IMC23_4294 when (BITSEL_u8_u1_4450_wire(0) /=  '0') else IMC22_4286;
    -- logger for split-operator MUX_4461_inst flow-through 
    process(IMD12_4462) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_4461_inst:flowthrough inputs: " & " BITSEL_u8_u1_4458_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4458_wire) & " IMC25_4310 = "& Convert_SLV_To_Hex_String(IMC25_4310) & " IMC24_4302 = "& Convert_SLV_To_Hex_String(IMC24_4302) & " outputs:" & " IMD12_4462= "  & Convert_SLV_To_Hex_String(IMD12_4462));
      --
    end process; 
    -- flow-through select operator MUX_4461_inst
    IMD12_4462 <= IMC25_4310 when (BITSEL_u8_u1_4458_wire(0) /=  '0') else IMC24_4302;
    -- logger for split-operator MUX_4469_inst flow-through 
    process(IMD13_4470) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_4469_inst:flowthrough inputs: " & " BITSEL_u8_u1_4466_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4466_wire) & " IMC27_4326 = "& Convert_SLV_To_Hex_String(IMC27_4326) & " IMC26_4318 = "& Convert_SLV_To_Hex_String(IMC26_4318) & " outputs:" & " IMD13_4470= "  & Convert_SLV_To_Hex_String(IMD13_4470));
      --
    end process; 
    -- flow-through select operator MUX_4469_inst
    IMD13_4470 <= IMC27_4326 when (BITSEL_u8_u1_4466_wire(0) /=  '0') else IMC26_4318;
    -- logger for split-operator MUX_4477_inst flow-through 
    process(IMD14_4478) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_4477_inst:flowthrough inputs: " & " BITSEL_u8_u1_4474_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4474_wire) & " IMC29_4342 = "& Convert_SLV_To_Hex_String(IMC29_4342) & " IMC28_4334 = "& Convert_SLV_To_Hex_String(IMC28_4334) & " outputs:" & " IMD14_4478= "  & Convert_SLV_To_Hex_String(IMD14_4478));
      --
    end process; 
    -- flow-through select operator MUX_4477_inst
    IMD14_4478 <= IMC29_4342 when (BITSEL_u8_u1_4474_wire(0) /=  '0') else IMC28_4334;
    -- logger for split-operator MUX_4485_inst flow-through 
    process(IMD15_4486) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_4485_inst:flowthrough inputs: " & " BITSEL_u8_u1_4482_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4482_wire) & " IMC31_4358 = "& Convert_SLV_To_Hex_String(IMC31_4358) & " IMC30_4350 = "& Convert_SLV_To_Hex_String(IMC30_4350) & " outputs:" & " IMD15_4486= "  & Convert_SLV_To_Hex_String(IMD15_4486));
      --
    end process; 
    -- flow-through select operator MUX_4485_inst
    IMD15_4486 <= IMC31_4358 when (BITSEL_u8_u1_4482_wire(0) /=  '0') else IMC30_4350;
    -- logger for split-operator MUX_4493_inst flow-through 
    process(IME0_4494) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_4493_inst:flowthrough inputs: " & " BITSEL_u8_u1_4490_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4490_wire) & " IMD1_4374 = "& Convert_SLV_To_Hex_String(IMD1_4374) & " IMD0_4366 = "& Convert_SLV_To_Hex_String(IMD0_4366) & " outputs:" & " IME0_4494= "  & Convert_SLV_To_Hex_String(IME0_4494));
      --
    end process; 
    -- flow-through select operator MUX_4493_inst
    IME0_4494 <= IMD1_4374 when (BITSEL_u8_u1_4490_wire(0) /=  '0') else IMD0_4366;
    -- logger for split-operator MUX_4501_inst flow-through 
    process(IME1_4502) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_4501_inst:flowthrough inputs: " & " BITSEL_u8_u1_4498_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4498_wire) & " IMD3_4390 = "& Convert_SLV_To_Hex_String(IMD3_4390) & " IMD2_4382 = "& Convert_SLV_To_Hex_String(IMD2_4382) & " outputs:" & " IME1_4502= "  & Convert_SLV_To_Hex_String(IME1_4502));
      --
    end process; 
    -- flow-through select operator MUX_4501_inst
    IME1_4502 <= IMD3_4390 when (BITSEL_u8_u1_4498_wire(0) /=  '0') else IMD2_4382;
    -- logger for split-operator MUX_4509_inst flow-through 
    process(IME2_4510) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_4509_inst:flowthrough inputs: " & " BITSEL_u8_u1_4506_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4506_wire) & " IMD5_4406 = "& Convert_SLV_To_Hex_String(IMD5_4406) & " IMD4_4398 = "& Convert_SLV_To_Hex_String(IMD4_4398) & " outputs:" & " IME2_4510= "  & Convert_SLV_To_Hex_String(IME2_4510));
      --
    end process; 
    -- flow-through select operator MUX_4509_inst
    IME2_4510 <= IMD5_4406 when (BITSEL_u8_u1_4506_wire(0) /=  '0') else IMD4_4398;
    -- logger for split-operator MUX_4517_inst flow-through 
    process(IME3_4518) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_4517_inst:flowthrough inputs: " & " BITSEL_u8_u1_4514_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4514_wire) & " IMD7_4422 = "& Convert_SLV_To_Hex_String(IMD7_4422) & " IMD6_4414 = "& Convert_SLV_To_Hex_String(IMD6_4414) & " outputs:" & " IME3_4518= "  & Convert_SLV_To_Hex_String(IME3_4518));
      --
    end process; 
    -- flow-through select operator MUX_4517_inst
    IME3_4518 <= IMD7_4422 when (BITSEL_u8_u1_4514_wire(0) /=  '0') else IMD6_4414;
    -- logger for split-operator MUX_4525_inst flow-through 
    process(IME4_4526) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_4525_inst:flowthrough inputs: " & " BITSEL_u8_u1_4522_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4522_wire) & " IMD9_4438 = "& Convert_SLV_To_Hex_String(IMD9_4438) & " IMD8_4430 = "& Convert_SLV_To_Hex_String(IMD8_4430) & " outputs:" & " IME4_4526= "  & Convert_SLV_To_Hex_String(IME4_4526));
      --
    end process; 
    -- flow-through select operator MUX_4525_inst
    IME4_4526 <= IMD9_4438 when (BITSEL_u8_u1_4522_wire(0) /=  '0') else IMD8_4430;
    -- logger for split-operator MUX_4533_inst flow-through 
    process(IME5_4534) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_4533_inst:flowthrough inputs: " & " BITSEL_u8_u1_4530_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4530_wire) & " IMD11_4454 = "& Convert_SLV_To_Hex_String(IMD11_4454) & " IMD10_4446 = "& Convert_SLV_To_Hex_String(IMD10_4446) & " outputs:" & " IME5_4534= "  & Convert_SLV_To_Hex_String(IME5_4534));
      --
    end process; 
    -- flow-through select operator MUX_4533_inst
    IME5_4534 <= IMD11_4454 when (BITSEL_u8_u1_4530_wire(0) /=  '0') else IMD10_4446;
    -- logger for split-operator MUX_4541_inst flow-through 
    process(IME6_4542) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_4541_inst:flowthrough inputs: " & " BITSEL_u8_u1_4538_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4538_wire) & " IMD13_4470 = "& Convert_SLV_To_Hex_String(IMD13_4470) & " IMD12_4462 = "& Convert_SLV_To_Hex_String(IMD12_4462) & " outputs:" & " IME6_4542= "  & Convert_SLV_To_Hex_String(IME6_4542));
      --
    end process; 
    -- flow-through select operator MUX_4541_inst
    IME6_4542 <= IMD13_4470 when (BITSEL_u8_u1_4538_wire(0) /=  '0') else IMD12_4462;
    -- logger for split-operator MUX_4549_inst flow-through 
    process(IME7_4550) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_4549_inst:flowthrough inputs: " & " BITSEL_u8_u1_4546_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4546_wire) & " IMD15_4486 = "& Convert_SLV_To_Hex_String(IMD15_4486) & " IMD14_4478 = "& Convert_SLV_To_Hex_String(IMD14_4478) & " outputs:" & " IME7_4550= "  & Convert_SLV_To_Hex_String(IME7_4550));
      --
    end process; 
    -- flow-through select operator MUX_4549_inst
    IME7_4550 <= IMD15_4486 when (BITSEL_u8_u1_4546_wire(0) /=  '0') else IMD14_4478;
    -- logger for split-operator MUX_4557_inst flow-through 
    process(IMF0_4558) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_4557_inst:flowthrough inputs: " & " BITSEL_u8_u1_4554_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4554_wire) & " IME1_4502 = "& Convert_SLV_To_Hex_String(IME1_4502) & " IME0_4494 = "& Convert_SLV_To_Hex_String(IME0_4494) & " outputs:" & " IMF0_4558= "  & Convert_SLV_To_Hex_String(IMF0_4558));
      --
    end process; 
    -- flow-through select operator MUX_4557_inst
    IMF0_4558 <= IME1_4502 when (BITSEL_u8_u1_4554_wire(0) /=  '0') else IME0_4494;
    -- logger for split-operator MUX_4565_inst flow-through 
    process(IMF1_4566) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_4565_inst:flowthrough inputs: " & " BITSEL_u8_u1_4562_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4562_wire) & " IME3_4518 = "& Convert_SLV_To_Hex_String(IME3_4518) & " IME2_4510 = "& Convert_SLV_To_Hex_String(IME2_4510) & " outputs:" & " IMF1_4566= "  & Convert_SLV_To_Hex_String(IMF1_4566));
      --
    end process; 
    -- flow-through select operator MUX_4565_inst
    IMF1_4566 <= IME3_4518 when (BITSEL_u8_u1_4562_wire(0) /=  '0') else IME2_4510;
    -- logger for split-operator MUX_4573_inst flow-through 
    process(IMF2_4574) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_4573_inst:flowthrough inputs: " & " BITSEL_u8_u1_4570_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4570_wire) & " IME5_4534 = "& Convert_SLV_To_Hex_String(IME5_4534) & " IME4_4526 = "& Convert_SLV_To_Hex_String(IME4_4526) & " outputs:" & " IMF2_4574= "  & Convert_SLV_To_Hex_String(IMF2_4574));
      --
    end process; 
    -- flow-through select operator MUX_4573_inst
    IMF2_4574 <= IME5_4534 when (BITSEL_u8_u1_4570_wire(0) /=  '0') else IME4_4526;
    -- logger for split-operator MUX_4581_inst flow-through 
    process(IMF3_4582) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_4581_inst:flowthrough inputs: " & " BITSEL_u8_u1_4578_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4578_wire) & " IME7_4550 = "& Convert_SLV_To_Hex_String(IME7_4550) & " IME6_4542 = "& Convert_SLV_To_Hex_String(IME6_4542) & " outputs:" & " IMF3_4582= "  & Convert_SLV_To_Hex_String(IMF3_4582));
      --
    end process; 
    -- flow-through select operator MUX_4581_inst
    IMF3_4582 <= IME7_4550 when (BITSEL_u8_u1_4578_wire(0) /=  '0') else IME6_4542;
    -- logger for split-operator MUX_4589_inst flow-through 
    process(IMG0_4590) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_4589_inst:flowthrough inputs: " & " BITSEL_u8_u1_4586_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4586_wire) & " IMF1_4566 = "& Convert_SLV_To_Hex_String(IMF1_4566) & " IMF0_4558 = "& Convert_SLV_To_Hex_String(IMF0_4558) & " outputs:" & " IMG0_4590= "  & Convert_SLV_To_Hex_String(IMG0_4590));
      --
    end process; 
    -- flow-through select operator MUX_4589_inst
    IMG0_4590 <= IMF1_4566 when (BITSEL_u8_u1_4586_wire(0) /=  '0') else IMF0_4558;
    -- logger for split-operator MUX_4597_inst flow-through 
    process(IMG1_4598) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_4597_inst:flowthrough inputs: " & " BITSEL_u8_u1_4594_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4594_wire) & " IMF3_4582 = "& Convert_SLV_To_Hex_String(IMF3_4582) & " IMF2_4574 = "& Convert_SLV_To_Hex_String(IMF2_4574) & " outputs:" & " IMG1_4598= "  & Convert_SLV_To_Hex_String(IMG1_4598));
      --
    end process; 
    -- flow-through select operator MUX_4597_inst
    IMG1_4598 <= IMF3_4582 when (BITSEL_u8_u1_4594_wire(0) /=  '0') else IMF2_4574;
    -- logger for split-operator MUX_4605_inst flow-through 
    process(s_out_buffer) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:MUX_4605_inst:flowthrough inputs: " & " BITSEL_u8_u1_4602_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4602_wire) & " IMG1_4598 = "& Convert_SLV_To_Hex_String(IMG1_4598) & " IMG0_4590 = "& Convert_SLV_To_Hex_String(IMG0_4590) & " outputs:" & " s_out_buffer= "  & Convert_SLV_To_Hex_String(s_out_buffer));
      --
    end process; 
    -- flow-through select operator MUX_4605_inst
    s_out_buffer <= IMG1_4598 when (BITSEL_u8_u1_4602_wire(0) /=  '0') else IMG0_4590;
    -- logger for split-operator BITSEL_u8_u1_2314_inst flow-through 
    process(BITSEL_u8_u1_2314_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_2314_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_2313_wire_constant = "& Convert_SLV_To_Hex_String(konst_2313_wire_constant) & " outputs:" & " BITSEL_u8_u1_2314_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_2314_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_2314_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2313_wire_constant, tmp_var);
      BITSEL_u8_u1_2314_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_2324_inst flow-through 
    process(BITSEL_u8_u1_2324_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_2324_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_2323_wire_constant = "& Convert_SLV_To_Hex_String(konst_2323_wire_constant) & " outputs:" & " BITSEL_u8_u1_2324_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_2324_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_2324_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2323_wire_constant, tmp_var);
      BITSEL_u8_u1_2324_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_2334_inst flow-through 
    process(BITSEL_u8_u1_2334_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_2334_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_2333_wire_constant = "& Convert_SLV_To_Hex_String(konst_2333_wire_constant) & " outputs:" & " BITSEL_u8_u1_2334_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_2334_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_2334_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2333_wire_constant, tmp_var);
      BITSEL_u8_u1_2334_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_2344_inst flow-through 
    process(BITSEL_u8_u1_2344_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_2344_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_2343_wire_constant = "& Convert_SLV_To_Hex_String(konst_2343_wire_constant) & " outputs:" & " BITSEL_u8_u1_2344_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_2344_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_2344_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2343_wire_constant, tmp_var);
      BITSEL_u8_u1_2344_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_2354_inst flow-through 
    process(BITSEL_u8_u1_2354_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_2354_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_2353_wire_constant = "& Convert_SLV_To_Hex_String(konst_2353_wire_constant) & " outputs:" & " BITSEL_u8_u1_2354_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_2354_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_2354_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2353_wire_constant, tmp_var);
      BITSEL_u8_u1_2354_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_2364_inst flow-through 
    process(BITSEL_u8_u1_2364_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_2364_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_2363_wire_constant = "& Convert_SLV_To_Hex_String(konst_2363_wire_constant) & " outputs:" & " BITSEL_u8_u1_2364_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_2364_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_2364_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2363_wire_constant, tmp_var);
      BITSEL_u8_u1_2364_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_2374_inst flow-through 
    process(BITSEL_u8_u1_2374_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_2374_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_2373_wire_constant = "& Convert_SLV_To_Hex_String(konst_2373_wire_constant) & " outputs:" & " BITSEL_u8_u1_2374_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_2374_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_2374_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2373_wire_constant, tmp_var);
      BITSEL_u8_u1_2374_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_2384_inst flow-through 
    process(BITSEL_u8_u1_2384_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_2384_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_2383_wire_constant = "& Convert_SLV_To_Hex_String(konst_2383_wire_constant) & " outputs:" & " BITSEL_u8_u1_2384_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_2384_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_2384_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2383_wire_constant, tmp_var);
      BITSEL_u8_u1_2384_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_2394_inst flow-through 
    process(BITSEL_u8_u1_2394_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_2394_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_2393_wire_constant = "& Convert_SLV_To_Hex_String(konst_2393_wire_constant) & " outputs:" & " BITSEL_u8_u1_2394_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_2394_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_2394_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2393_wire_constant, tmp_var);
      BITSEL_u8_u1_2394_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_2404_inst flow-through 
    process(BITSEL_u8_u1_2404_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_2404_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_2403_wire_constant = "& Convert_SLV_To_Hex_String(konst_2403_wire_constant) & " outputs:" & " BITSEL_u8_u1_2404_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_2404_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_2404_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2403_wire_constant, tmp_var);
      BITSEL_u8_u1_2404_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_2414_inst flow-through 
    process(BITSEL_u8_u1_2414_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_2414_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_2413_wire_constant = "& Convert_SLV_To_Hex_String(konst_2413_wire_constant) & " outputs:" & " BITSEL_u8_u1_2414_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_2414_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_2414_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2413_wire_constant, tmp_var);
      BITSEL_u8_u1_2414_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_2424_inst flow-through 
    process(BITSEL_u8_u1_2424_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_2424_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_2423_wire_constant = "& Convert_SLV_To_Hex_String(konst_2423_wire_constant) & " outputs:" & " BITSEL_u8_u1_2424_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_2424_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_2424_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2423_wire_constant, tmp_var);
      BITSEL_u8_u1_2424_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_2434_inst flow-through 
    process(BITSEL_u8_u1_2434_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_2434_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_2433_wire_constant = "& Convert_SLV_To_Hex_String(konst_2433_wire_constant) & " outputs:" & " BITSEL_u8_u1_2434_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_2434_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_2434_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2433_wire_constant, tmp_var);
      BITSEL_u8_u1_2434_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_2444_inst flow-through 
    process(BITSEL_u8_u1_2444_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_2444_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_2443_wire_constant = "& Convert_SLV_To_Hex_String(konst_2443_wire_constant) & " outputs:" & " BITSEL_u8_u1_2444_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_2444_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_2444_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2443_wire_constant, tmp_var);
      BITSEL_u8_u1_2444_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_2454_inst flow-through 
    process(BITSEL_u8_u1_2454_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_2454_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_2453_wire_constant = "& Convert_SLV_To_Hex_String(konst_2453_wire_constant) & " outputs:" & " BITSEL_u8_u1_2454_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_2454_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_2454_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2453_wire_constant, tmp_var);
      BITSEL_u8_u1_2454_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_2464_inst flow-through 
    process(BITSEL_u8_u1_2464_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_2464_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_2463_wire_constant = "& Convert_SLV_To_Hex_String(konst_2463_wire_constant) & " outputs:" & " BITSEL_u8_u1_2464_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_2464_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_2464_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2463_wire_constant, tmp_var);
      BITSEL_u8_u1_2464_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_2474_inst flow-through 
    process(BITSEL_u8_u1_2474_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_2474_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_2473_wire_constant = "& Convert_SLV_To_Hex_String(konst_2473_wire_constant) & " outputs:" & " BITSEL_u8_u1_2474_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_2474_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_2474_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2473_wire_constant, tmp_var);
      BITSEL_u8_u1_2474_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_2484_inst flow-through 
    process(BITSEL_u8_u1_2484_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_2484_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_2483_wire_constant = "& Convert_SLV_To_Hex_String(konst_2483_wire_constant) & " outputs:" & " BITSEL_u8_u1_2484_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_2484_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_2484_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2483_wire_constant, tmp_var);
      BITSEL_u8_u1_2484_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_2494_inst flow-through 
    process(BITSEL_u8_u1_2494_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_2494_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_2493_wire_constant = "& Convert_SLV_To_Hex_String(konst_2493_wire_constant) & " outputs:" & " BITSEL_u8_u1_2494_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_2494_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_2494_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2493_wire_constant, tmp_var);
      BITSEL_u8_u1_2494_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_2504_inst flow-through 
    process(BITSEL_u8_u1_2504_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_2504_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_2503_wire_constant = "& Convert_SLV_To_Hex_String(konst_2503_wire_constant) & " outputs:" & " BITSEL_u8_u1_2504_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_2504_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_2504_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2503_wire_constant, tmp_var);
      BITSEL_u8_u1_2504_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_2514_inst flow-through 
    process(BITSEL_u8_u1_2514_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_2514_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_2513_wire_constant = "& Convert_SLV_To_Hex_String(konst_2513_wire_constant) & " outputs:" & " BITSEL_u8_u1_2514_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_2514_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_2514_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2513_wire_constant, tmp_var);
      BITSEL_u8_u1_2514_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_2524_inst flow-through 
    process(BITSEL_u8_u1_2524_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_2524_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_2523_wire_constant = "& Convert_SLV_To_Hex_String(konst_2523_wire_constant) & " outputs:" & " BITSEL_u8_u1_2524_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_2524_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_2524_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2523_wire_constant, tmp_var);
      BITSEL_u8_u1_2524_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_2534_inst flow-through 
    process(BITSEL_u8_u1_2534_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_2534_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_2533_wire_constant = "& Convert_SLV_To_Hex_String(konst_2533_wire_constant) & " outputs:" & " BITSEL_u8_u1_2534_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_2534_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_2534_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2533_wire_constant, tmp_var);
      BITSEL_u8_u1_2534_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_2544_inst flow-through 
    process(BITSEL_u8_u1_2544_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_2544_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_2543_wire_constant = "& Convert_SLV_To_Hex_String(konst_2543_wire_constant) & " outputs:" & " BITSEL_u8_u1_2544_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_2544_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_2544_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2543_wire_constant, tmp_var);
      BITSEL_u8_u1_2544_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_2554_inst flow-through 
    process(BITSEL_u8_u1_2554_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_2554_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_2553_wire_constant = "& Convert_SLV_To_Hex_String(konst_2553_wire_constant) & " outputs:" & " BITSEL_u8_u1_2554_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_2554_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_2554_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2553_wire_constant, tmp_var);
      BITSEL_u8_u1_2554_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_2564_inst flow-through 
    process(BITSEL_u8_u1_2564_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_2564_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_2563_wire_constant = "& Convert_SLV_To_Hex_String(konst_2563_wire_constant) & " outputs:" & " BITSEL_u8_u1_2564_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_2564_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_2564_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2563_wire_constant, tmp_var);
      BITSEL_u8_u1_2564_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_2574_inst flow-through 
    process(BITSEL_u8_u1_2574_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_2574_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_2573_wire_constant = "& Convert_SLV_To_Hex_String(konst_2573_wire_constant) & " outputs:" & " BITSEL_u8_u1_2574_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_2574_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_2574_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2573_wire_constant, tmp_var);
      BITSEL_u8_u1_2574_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_2584_inst flow-through 
    process(BITSEL_u8_u1_2584_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_2584_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_2583_wire_constant = "& Convert_SLV_To_Hex_String(konst_2583_wire_constant) & " outputs:" & " BITSEL_u8_u1_2584_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_2584_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_2584_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2583_wire_constant, tmp_var);
      BITSEL_u8_u1_2584_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_2594_inst flow-through 
    process(BITSEL_u8_u1_2594_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_2594_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_2593_wire_constant = "& Convert_SLV_To_Hex_String(konst_2593_wire_constant) & " outputs:" & " BITSEL_u8_u1_2594_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_2594_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_2594_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2593_wire_constant, tmp_var);
      BITSEL_u8_u1_2594_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_2604_inst flow-through 
    process(BITSEL_u8_u1_2604_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_2604_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_2603_wire_constant = "& Convert_SLV_To_Hex_String(konst_2603_wire_constant) & " outputs:" & " BITSEL_u8_u1_2604_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_2604_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_2604_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2603_wire_constant, tmp_var);
      BITSEL_u8_u1_2604_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_2614_inst flow-through 
    process(BITSEL_u8_u1_2614_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_2614_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_2613_wire_constant = "& Convert_SLV_To_Hex_String(konst_2613_wire_constant) & " outputs:" & " BITSEL_u8_u1_2614_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_2614_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_2614_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2613_wire_constant, tmp_var);
      BITSEL_u8_u1_2614_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_2624_inst flow-through 
    process(BITSEL_u8_u1_2624_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_2624_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_2623_wire_constant = "& Convert_SLV_To_Hex_String(konst_2623_wire_constant) & " outputs:" & " BITSEL_u8_u1_2624_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_2624_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_2624_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2623_wire_constant, tmp_var);
      BITSEL_u8_u1_2624_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_2634_inst flow-through 
    process(BITSEL_u8_u1_2634_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_2634_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_2633_wire_constant = "& Convert_SLV_To_Hex_String(konst_2633_wire_constant) & " outputs:" & " BITSEL_u8_u1_2634_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_2634_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_2634_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2633_wire_constant, tmp_var);
      BITSEL_u8_u1_2634_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_2644_inst flow-through 
    process(BITSEL_u8_u1_2644_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_2644_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_2643_wire_constant = "& Convert_SLV_To_Hex_String(konst_2643_wire_constant) & " outputs:" & " BITSEL_u8_u1_2644_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_2644_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_2644_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2643_wire_constant, tmp_var);
      BITSEL_u8_u1_2644_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_2654_inst flow-through 
    process(BITSEL_u8_u1_2654_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_2654_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_2653_wire_constant = "& Convert_SLV_To_Hex_String(konst_2653_wire_constant) & " outputs:" & " BITSEL_u8_u1_2654_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_2654_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_2654_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2653_wire_constant, tmp_var);
      BITSEL_u8_u1_2654_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_2664_inst flow-through 
    process(BITSEL_u8_u1_2664_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_2664_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_2663_wire_constant = "& Convert_SLV_To_Hex_String(konst_2663_wire_constant) & " outputs:" & " BITSEL_u8_u1_2664_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_2664_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_2664_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2663_wire_constant, tmp_var);
      BITSEL_u8_u1_2664_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_2674_inst flow-through 
    process(BITSEL_u8_u1_2674_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_2674_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_2673_wire_constant = "& Convert_SLV_To_Hex_String(konst_2673_wire_constant) & " outputs:" & " BITSEL_u8_u1_2674_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_2674_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_2674_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2673_wire_constant, tmp_var);
      BITSEL_u8_u1_2674_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_2684_inst flow-through 
    process(BITSEL_u8_u1_2684_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_2684_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_2683_wire_constant = "& Convert_SLV_To_Hex_String(konst_2683_wire_constant) & " outputs:" & " BITSEL_u8_u1_2684_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_2684_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_2684_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2683_wire_constant, tmp_var);
      BITSEL_u8_u1_2684_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_2694_inst flow-through 
    process(BITSEL_u8_u1_2694_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_2694_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_2693_wire_constant = "& Convert_SLV_To_Hex_String(konst_2693_wire_constant) & " outputs:" & " BITSEL_u8_u1_2694_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_2694_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_2694_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2693_wire_constant, tmp_var);
      BITSEL_u8_u1_2694_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_2704_inst flow-through 
    process(BITSEL_u8_u1_2704_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_2704_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_2703_wire_constant = "& Convert_SLV_To_Hex_String(konst_2703_wire_constant) & " outputs:" & " BITSEL_u8_u1_2704_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_2704_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_2704_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2703_wire_constant, tmp_var);
      BITSEL_u8_u1_2704_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_2714_inst flow-through 
    process(BITSEL_u8_u1_2714_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_2714_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_2713_wire_constant = "& Convert_SLV_To_Hex_String(konst_2713_wire_constant) & " outputs:" & " BITSEL_u8_u1_2714_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_2714_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_2714_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2713_wire_constant, tmp_var);
      BITSEL_u8_u1_2714_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_2724_inst flow-through 
    process(BITSEL_u8_u1_2724_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_2724_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_2723_wire_constant = "& Convert_SLV_To_Hex_String(konst_2723_wire_constant) & " outputs:" & " BITSEL_u8_u1_2724_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_2724_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_2724_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2723_wire_constant, tmp_var);
      BITSEL_u8_u1_2724_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_2734_inst flow-through 
    process(BITSEL_u8_u1_2734_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_2734_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_2733_wire_constant = "& Convert_SLV_To_Hex_String(konst_2733_wire_constant) & " outputs:" & " BITSEL_u8_u1_2734_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_2734_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_2734_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2733_wire_constant, tmp_var);
      BITSEL_u8_u1_2734_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_2744_inst flow-through 
    process(BITSEL_u8_u1_2744_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_2744_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_2743_wire_constant = "& Convert_SLV_To_Hex_String(konst_2743_wire_constant) & " outputs:" & " BITSEL_u8_u1_2744_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_2744_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_2744_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2743_wire_constant, tmp_var);
      BITSEL_u8_u1_2744_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_2754_inst flow-through 
    process(BITSEL_u8_u1_2754_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_2754_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_2753_wire_constant = "& Convert_SLV_To_Hex_String(konst_2753_wire_constant) & " outputs:" & " BITSEL_u8_u1_2754_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_2754_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_2754_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2753_wire_constant, tmp_var);
      BITSEL_u8_u1_2754_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_2764_inst flow-through 
    process(BITSEL_u8_u1_2764_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_2764_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_2763_wire_constant = "& Convert_SLV_To_Hex_String(konst_2763_wire_constant) & " outputs:" & " BITSEL_u8_u1_2764_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_2764_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_2764_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2763_wire_constant, tmp_var);
      BITSEL_u8_u1_2764_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_2774_inst flow-through 
    process(BITSEL_u8_u1_2774_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_2774_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_2773_wire_constant = "& Convert_SLV_To_Hex_String(konst_2773_wire_constant) & " outputs:" & " BITSEL_u8_u1_2774_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_2774_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_2774_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2773_wire_constant, tmp_var);
      BITSEL_u8_u1_2774_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_2784_inst flow-through 
    process(BITSEL_u8_u1_2784_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_2784_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_2783_wire_constant = "& Convert_SLV_To_Hex_String(konst_2783_wire_constant) & " outputs:" & " BITSEL_u8_u1_2784_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_2784_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_2784_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2783_wire_constant, tmp_var);
      BITSEL_u8_u1_2784_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_2794_inst flow-through 
    process(BITSEL_u8_u1_2794_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_2794_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_2793_wire_constant = "& Convert_SLV_To_Hex_String(konst_2793_wire_constant) & " outputs:" & " BITSEL_u8_u1_2794_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_2794_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_2794_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2793_wire_constant, tmp_var);
      BITSEL_u8_u1_2794_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_2804_inst flow-through 
    process(BITSEL_u8_u1_2804_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_2804_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_2803_wire_constant = "& Convert_SLV_To_Hex_String(konst_2803_wire_constant) & " outputs:" & " BITSEL_u8_u1_2804_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_2804_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_2804_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2803_wire_constant, tmp_var);
      BITSEL_u8_u1_2804_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_2814_inst flow-through 
    process(BITSEL_u8_u1_2814_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_2814_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_2813_wire_constant = "& Convert_SLV_To_Hex_String(konst_2813_wire_constant) & " outputs:" & " BITSEL_u8_u1_2814_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_2814_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_2814_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2813_wire_constant, tmp_var);
      BITSEL_u8_u1_2814_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_2824_inst flow-through 
    process(BITSEL_u8_u1_2824_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_2824_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_2823_wire_constant = "& Convert_SLV_To_Hex_String(konst_2823_wire_constant) & " outputs:" & " BITSEL_u8_u1_2824_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_2824_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_2824_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2823_wire_constant, tmp_var);
      BITSEL_u8_u1_2824_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_2834_inst flow-through 
    process(BITSEL_u8_u1_2834_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_2834_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_2833_wire_constant = "& Convert_SLV_To_Hex_String(konst_2833_wire_constant) & " outputs:" & " BITSEL_u8_u1_2834_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_2834_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_2834_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2833_wire_constant, tmp_var);
      BITSEL_u8_u1_2834_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_2844_inst flow-through 
    process(BITSEL_u8_u1_2844_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_2844_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_2843_wire_constant = "& Convert_SLV_To_Hex_String(konst_2843_wire_constant) & " outputs:" & " BITSEL_u8_u1_2844_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_2844_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_2844_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2843_wire_constant, tmp_var);
      BITSEL_u8_u1_2844_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_2854_inst flow-through 
    process(BITSEL_u8_u1_2854_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_2854_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_2853_wire_constant = "& Convert_SLV_To_Hex_String(konst_2853_wire_constant) & " outputs:" & " BITSEL_u8_u1_2854_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_2854_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_2854_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2853_wire_constant, tmp_var);
      BITSEL_u8_u1_2854_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_2864_inst flow-through 
    process(BITSEL_u8_u1_2864_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_2864_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_2863_wire_constant = "& Convert_SLV_To_Hex_String(konst_2863_wire_constant) & " outputs:" & " BITSEL_u8_u1_2864_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_2864_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_2864_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2863_wire_constant, tmp_var);
      BITSEL_u8_u1_2864_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_2874_inst flow-through 
    process(BITSEL_u8_u1_2874_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_2874_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_2873_wire_constant = "& Convert_SLV_To_Hex_String(konst_2873_wire_constant) & " outputs:" & " BITSEL_u8_u1_2874_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_2874_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_2874_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2873_wire_constant, tmp_var);
      BITSEL_u8_u1_2874_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_2884_inst flow-through 
    process(BITSEL_u8_u1_2884_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_2884_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_2883_wire_constant = "& Convert_SLV_To_Hex_String(konst_2883_wire_constant) & " outputs:" & " BITSEL_u8_u1_2884_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_2884_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_2884_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2883_wire_constant, tmp_var);
      BITSEL_u8_u1_2884_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_2894_inst flow-through 
    process(BITSEL_u8_u1_2894_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_2894_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_2893_wire_constant = "& Convert_SLV_To_Hex_String(konst_2893_wire_constant) & " outputs:" & " BITSEL_u8_u1_2894_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_2894_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_2894_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2893_wire_constant, tmp_var);
      BITSEL_u8_u1_2894_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_2904_inst flow-through 
    process(BITSEL_u8_u1_2904_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_2904_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_2903_wire_constant = "& Convert_SLV_To_Hex_String(konst_2903_wire_constant) & " outputs:" & " BITSEL_u8_u1_2904_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_2904_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_2904_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2903_wire_constant, tmp_var);
      BITSEL_u8_u1_2904_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_2914_inst flow-through 
    process(BITSEL_u8_u1_2914_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_2914_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_2913_wire_constant = "& Convert_SLV_To_Hex_String(konst_2913_wire_constant) & " outputs:" & " BITSEL_u8_u1_2914_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_2914_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_2914_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2913_wire_constant, tmp_var);
      BITSEL_u8_u1_2914_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_2924_inst flow-through 
    process(BITSEL_u8_u1_2924_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_2924_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_2923_wire_constant = "& Convert_SLV_To_Hex_String(konst_2923_wire_constant) & " outputs:" & " BITSEL_u8_u1_2924_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_2924_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_2924_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2923_wire_constant, tmp_var);
      BITSEL_u8_u1_2924_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_2934_inst flow-through 
    process(BITSEL_u8_u1_2934_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_2934_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_2933_wire_constant = "& Convert_SLV_To_Hex_String(konst_2933_wire_constant) & " outputs:" & " BITSEL_u8_u1_2934_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_2934_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_2934_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2933_wire_constant, tmp_var);
      BITSEL_u8_u1_2934_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_2944_inst flow-through 
    process(BITSEL_u8_u1_2944_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_2944_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_2943_wire_constant = "& Convert_SLV_To_Hex_String(konst_2943_wire_constant) & " outputs:" & " BITSEL_u8_u1_2944_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_2944_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_2944_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2943_wire_constant, tmp_var);
      BITSEL_u8_u1_2944_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_2954_inst flow-through 
    process(BITSEL_u8_u1_2954_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_2954_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_2953_wire_constant = "& Convert_SLV_To_Hex_String(konst_2953_wire_constant) & " outputs:" & " BITSEL_u8_u1_2954_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_2954_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_2954_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2953_wire_constant, tmp_var);
      BITSEL_u8_u1_2954_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_2964_inst flow-through 
    process(BITSEL_u8_u1_2964_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_2964_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_2963_wire_constant = "& Convert_SLV_To_Hex_String(konst_2963_wire_constant) & " outputs:" & " BITSEL_u8_u1_2964_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_2964_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_2964_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2963_wire_constant, tmp_var);
      BITSEL_u8_u1_2964_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_2974_inst flow-through 
    process(BITSEL_u8_u1_2974_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_2974_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_2973_wire_constant = "& Convert_SLV_To_Hex_String(konst_2973_wire_constant) & " outputs:" & " BITSEL_u8_u1_2974_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_2974_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_2974_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2973_wire_constant, tmp_var);
      BITSEL_u8_u1_2974_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_2984_inst flow-through 
    process(BITSEL_u8_u1_2984_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_2984_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_2983_wire_constant = "& Convert_SLV_To_Hex_String(konst_2983_wire_constant) & " outputs:" & " BITSEL_u8_u1_2984_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_2984_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_2984_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2983_wire_constant, tmp_var);
      BITSEL_u8_u1_2984_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_2994_inst flow-through 
    process(BITSEL_u8_u1_2994_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_2994_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_2993_wire_constant = "& Convert_SLV_To_Hex_String(konst_2993_wire_constant) & " outputs:" & " BITSEL_u8_u1_2994_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_2994_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_2994_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2993_wire_constant, tmp_var);
      BITSEL_u8_u1_2994_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3004_inst flow-through 
    process(BITSEL_u8_u1_3004_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3004_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3003_wire_constant = "& Convert_SLV_To_Hex_String(konst_3003_wire_constant) & " outputs:" & " BITSEL_u8_u1_3004_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3004_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3004_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3003_wire_constant, tmp_var);
      BITSEL_u8_u1_3004_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3014_inst flow-through 
    process(BITSEL_u8_u1_3014_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3014_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3013_wire_constant = "& Convert_SLV_To_Hex_String(konst_3013_wire_constant) & " outputs:" & " BITSEL_u8_u1_3014_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3014_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3014_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3013_wire_constant, tmp_var);
      BITSEL_u8_u1_3014_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3024_inst flow-through 
    process(BITSEL_u8_u1_3024_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3024_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3023_wire_constant = "& Convert_SLV_To_Hex_String(konst_3023_wire_constant) & " outputs:" & " BITSEL_u8_u1_3024_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3024_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3024_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3023_wire_constant, tmp_var);
      BITSEL_u8_u1_3024_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3034_inst flow-through 
    process(BITSEL_u8_u1_3034_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3034_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3033_wire_constant = "& Convert_SLV_To_Hex_String(konst_3033_wire_constant) & " outputs:" & " BITSEL_u8_u1_3034_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3034_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3034_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3033_wire_constant, tmp_var);
      BITSEL_u8_u1_3034_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3044_inst flow-through 
    process(BITSEL_u8_u1_3044_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3044_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3043_wire_constant = "& Convert_SLV_To_Hex_String(konst_3043_wire_constant) & " outputs:" & " BITSEL_u8_u1_3044_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3044_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3044_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3043_wire_constant, tmp_var);
      BITSEL_u8_u1_3044_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3054_inst flow-through 
    process(BITSEL_u8_u1_3054_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3054_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3053_wire_constant = "& Convert_SLV_To_Hex_String(konst_3053_wire_constant) & " outputs:" & " BITSEL_u8_u1_3054_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3054_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3054_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3053_wire_constant, tmp_var);
      BITSEL_u8_u1_3054_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3064_inst flow-through 
    process(BITSEL_u8_u1_3064_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3064_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3063_wire_constant = "& Convert_SLV_To_Hex_String(konst_3063_wire_constant) & " outputs:" & " BITSEL_u8_u1_3064_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3064_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3064_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3063_wire_constant, tmp_var);
      BITSEL_u8_u1_3064_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3074_inst flow-through 
    process(BITSEL_u8_u1_3074_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3074_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3073_wire_constant = "& Convert_SLV_To_Hex_String(konst_3073_wire_constant) & " outputs:" & " BITSEL_u8_u1_3074_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3074_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3074_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3073_wire_constant, tmp_var);
      BITSEL_u8_u1_3074_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3084_inst flow-through 
    process(BITSEL_u8_u1_3084_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3084_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3083_wire_constant = "& Convert_SLV_To_Hex_String(konst_3083_wire_constant) & " outputs:" & " BITSEL_u8_u1_3084_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3084_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3084_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3083_wire_constant, tmp_var);
      BITSEL_u8_u1_3084_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3094_inst flow-through 
    process(BITSEL_u8_u1_3094_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3094_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3093_wire_constant = "& Convert_SLV_To_Hex_String(konst_3093_wire_constant) & " outputs:" & " BITSEL_u8_u1_3094_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3094_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3094_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3093_wire_constant, tmp_var);
      BITSEL_u8_u1_3094_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3104_inst flow-through 
    process(BITSEL_u8_u1_3104_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3104_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3103_wire_constant = "& Convert_SLV_To_Hex_String(konst_3103_wire_constant) & " outputs:" & " BITSEL_u8_u1_3104_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3104_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3104_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3103_wire_constant, tmp_var);
      BITSEL_u8_u1_3104_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3114_inst flow-through 
    process(BITSEL_u8_u1_3114_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3114_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3113_wire_constant = "& Convert_SLV_To_Hex_String(konst_3113_wire_constant) & " outputs:" & " BITSEL_u8_u1_3114_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3114_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3114_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3113_wire_constant, tmp_var);
      BITSEL_u8_u1_3114_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3124_inst flow-through 
    process(BITSEL_u8_u1_3124_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3124_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3123_wire_constant = "& Convert_SLV_To_Hex_String(konst_3123_wire_constant) & " outputs:" & " BITSEL_u8_u1_3124_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3124_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3124_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3123_wire_constant, tmp_var);
      BITSEL_u8_u1_3124_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3134_inst flow-through 
    process(BITSEL_u8_u1_3134_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3134_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3133_wire_constant = "& Convert_SLV_To_Hex_String(konst_3133_wire_constant) & " outputs:" & " BITSEL_u8_u1_3134_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3134_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3134_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3133_wire_constant, tmp_var);
      BITSEL_u8_u1_3134_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3144_inst flow-through 
    process(BITSEL_u8_u1_3144_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3144_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3143_wire_constant = "& Convert_SLV_To_Hex_String(konst_3143_wire_constant) & " outputs:" & " BITSEL_u8_u1_3144_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3144_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3144_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3143_wire_constant, tmp_var);
      BITSEL_u8_u1_3144_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3154_inst flow-through 
    process(BITSEL_u8_u1_3154_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3154_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3153_wire_constant = "& Convert_SLV_To_Hex_String(konst_3153_wire_constant) & " outputs:" & " BITSEL_u8_u1_3154_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3154_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3154_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3153_wire_constant, tmp_var);
      BITSEL_u8_u1_3154_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3164_inst flow-through 
    process(BITSEL_u8_u1_3164_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3164_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3163_wire_constant = "& Convert_SLV_To_Hex_String(konst_3163_wire_constant) & " outputs:" & " BITSEL_u8_u1_3164_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3164_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3164_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3163_wire_constant, tmp_var);
      BITSEL_u8_u1_3164_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3174_inst flow-through 
    process(BITSEL_u8_u1_3174_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3174_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3173_wire_constant = "& Convert_SLV_To_Hex_String(konst_3173_wire_constant) & " outputs:" & " BITSEL_u8_u1_3174_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3174_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3174_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3173_wire_constant, tmp_var);
      BITSEL_u8_u1_3174_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3184_inst flow-through 
    process(BITSEL_u8_u1_3184_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3184_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3183_wire_constant = "& Convert_SLV_To_Hex_String(konst_3183_wire_constant) & " outputs:" & " BITSEL_u8_u1_3184_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3184_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3184_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3183_wire_constant, tmp_var);
      BITSEL_u8_u1_3184_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3194_inst flow-through 
    process(BITSEL_u8_u1_3194_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3194_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3193_wire_constant = "& Convert_SLV_To_Hex_String(konst_3193_wire_constant) & " outputs:" & " BITSEL_u8_u1_3194_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3194_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3194_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3193_wire_constant, tmp_var);
      BITSEL_u8_u1_3194_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3204_inst flow-through 
    process(BITSEL_u8_u1_3204_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3204_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3203_wire_constant = "& Convert_SLV_To_Hex_String(konst_3203_wire_constant) & " outputs:" & " BITSEL_u8_u1_3204_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3204_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3204_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3203_wire_constant, tmp_var);
      BITSEL_u8_u1_3204_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3214_inst flow-through 
    process(BITSEL_u8_u1_3214_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3214_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3213_wire_constant = "& Convert_SLV_To_Hex_String(konst_3213_wire_constant) & " outputs:" & " BITSEL_u8_u1_3214_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3214_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3214_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3213_wire_constant, tmp_var);
      BITSEL_u8_u1_3214_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3224_inst flow-through 
    process(BITSEL_u8_u1_3224_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3224_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3223_wire_constant = "& Convert_SLV_To_Hex_String(konst_3223_wire_constant) & " outputs:" & " BITSEL_u8_u1_3224_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3224_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3224_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3223_wire_constant, tmp_var);
      BITSEL_u8_u1_3224_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3234_inst flow-through 
    process(BITSEL_u8_u1_3234_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3234_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3233_wire_constant = "& Convert_SLV_To_Hex_String(konst_3233_wire_constant) & " outputs:" & " BITSEL_u8_u1_3234_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3234_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3234_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3233_wire_constant, tmp_var);
      BITSEL_u8_u1_3234_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3244_inst flow-through 
    process(BITSEL_u8_u1_3244_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3244_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3243_wire_constant = "& Convert_SLV_To_Hex_String(konst_3243_wire_constant) & " outputs:" & " BITSEL_u8_u1_3244_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3244_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3244_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3243_wire_constant, tmp_var);
      BITSEL_u8_u1_3244_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3254_inst flow-through 
    process(BITSEL_u8_u1_3254_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3254_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3253_wire_constant = "& Convert_SLV_To_Hex_String(konst_3253_wire_constant) & " outputs:" & " BITSEL_u8_u1_3254_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3254_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3254_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3253_wire_constant, tmp_var);
      BITSEL_u8_u1_3254_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3264_inst flow-through 
    process(BITSEL_u8_u1_3264_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3264_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3263_wire_constant = "& Convert_SLV_To_Hex_String(konst_3263_wire_constant) & " outputs:" & " BITSEL_u8_u1_3264_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3264_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3264_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3263_wire_constant, tmp_var);
      BITSEL_u8_u1_3264_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3274_inst flow-through 
    process(BITSEL_u8_u1_3274_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3274_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3273_wire_constant = "& Convert_SLV_To_Hex_String(konst_3273_wire_constant) & " outputs:" & " BITSEL_u8_u1_3274_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3274_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3274_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3273_wire_constant, tmp_var);
      BITSEL_u8_u1_3274_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3284_inst flow-through 
    process(BITSEL_u8_u1_3284_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3284_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3283_wire_constant = "& Convert_SLV_To_Hex_String(konst_3283_wire_constant) & " outputs:" & " BITSEL_u8_u1_3284_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3284_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3284_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3283_wire_constant, tmp_var);
      BITSEL_u8_u1_3284_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3294_inst flow-through 
    process(BITSEL_u8_u1_3294_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3294_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3293_wire_constant = "& Convert_SLV_To_Hex_String(konst_3293_wire_constant) & " outputs:" & " BITSEL_u8_u1_3294_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3294_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3294_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3293_wire_constant, tmp_var);
      BITSEL_u8_u1_3294_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3304_inst flow-through 
    process(BITSEL_u8_u1_3304_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3304_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3303_wire_constant = "& Convert_SLV_To_Hex_String(konst_3303_wire_constant) & " outputs:" & " BITSEL_u8_u1_3304_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3304_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3304_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3303_wire_constant, tmp_var);
      BITSEL_u8_u1_3304_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3314_inst flow-through 
    process(BITSEL_u8_u1_3314_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3314_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3313_wire_constant = "& Convert_SLV_To_Hex_String(konst_3313_wire_constant) & " outputs:" & " BITSEL_u8_u1_3314_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3314_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3314_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3313_wire_constant, tmp_var);
      BITSEL_u8_u1_3314_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3324_inst flow-through 
    process(BITSEL_u8_u1_3324_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3324_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3323_wire_constant = "& Convert_SLV_To_Hex_String(konst_3323_wire_constant) & " outputs:" & " BITSEL_u8_u1_3324_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3324_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3324_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3323_wire_constant, tmp_var);
      BITSEL_u8_u1_3324_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3334_inst flow-through 
    process(BITSEL_u8_u1_3334_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3334_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3333_wire_constant = "& Convert_SLV_To_Hex_String(konst_3333_wire_constant) & " outputs:" & " BITSEL_u8_u1_3334_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3334_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3334_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3333_wire_constant, tmp_var);
      BITSEL_u8_u1_3334_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3344_inst flow-through 
    process(BITSEL_u8_u1_3344_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3344_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3343_wire_constant = "& Convert_SLV_To_Hex_String(konst_3343_wire_constant) & " outputs:" & " BITSEL_u8_u1_3344_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3344_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3344_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3343_wire_constant, tmp_var);
      BITSEL_u8_u1_3344_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3354_inst flow-through 
    process(BITSEL_u8_u1_3354_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3354_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3353_wire_constant = "& Convert_SLV_To_Hex_String(konst_3353_wire_constant) & " outputs:" & " BITSEL_u8_u1_3354_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3354_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3354_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3353_wire_constant, tmp_var);
      BITSEL_u8_u1_3354_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3364_inst flow-through 
    process(BITSEL_u8_u1_3364_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3364_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3363_wire_constant = "& Convert_SLV_To_Hex_String(konst_3363_wire_constant) & " outputs:" & " BITSEL_u8_u1_3364_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3364_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3364_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3363_wire_constant, tmp_var);
      BITSEL_u8_u1_3364_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3374_inst flow-through 
    process(BITSEL_u8_u1_3374_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3374_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3373_wire_constant = "& Convert_SLV_To_Hex_String(konst_3373_wire_constant) & " outputs:" & " BITSEL_u8_u1_3374_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3374_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3374_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3373_wire_constant, tmp_var);
      BITSEL_u8_u1_3374_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3384_inst flow-through 
    process(BITSEL_u8_u1_3384_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3384_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3383_wire_constant = "& Convert_SLV_To_Hex_String(konst_3383_wire_constant) & " outputs:" & " BITSEL_u8_u1_3384_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3384_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3384_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3383_wire_constant, tmp_var);
      BITSEL_u8_u1_3384_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3394_inst flow-through 
    process(BITSEL_u8_u1_3394_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3394_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3393_wire_constant = "& Convert_SLV_To_Hex_String(konst_3393_wire_constant) & " outputs:" & " BITSEL_u8_u1_3394_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3394_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3394_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3393_wire_constant, tmp_var);
      BITSEL_u8_u1_3394_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3404_inst flow-through 
    process(BITSEL_u8_u1_3404_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3404_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3403_wire_constant = "& Convert_SLV_To_Hex_String(konst_3403_wire_constant) & " outputs:" & " BITSEL_u8_u1_3404_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3404_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3404_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3403_wire_constant, tmp_var);
      BITSEL_u8_u1_3404_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3414_inst flow-through 
    process(BITSEL_u8_u1_3414_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3414_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3413_wire_constant = "& Convert_SLV_To_Hex_String(konst_3413_wire_constant) & " outputs:" & " BITSEL_u8_u1_3414_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3414_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3414_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3413_wire_constant, tmp_var);
      BITSEL_u8_u1_3414_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3424_inst flow-through 
    process(BITSEL_u8_u1_3424_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3424_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3423_wire_constant = "& Convert_SLV_To_Hex_String(konst_3423_wire_constant) & " outputs:" & " BITSEL_u8_u1_3424_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3424_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3424_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3423_wire_constant, tmp_var);
      BITSEL_u8_u1_3424_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3434_inst flow-through 
    process(BITSEL_u8_u1_3434_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3434_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3433_wire_constant = "& Convert_SLV_To_Hex_String(konst_3433_wire_constant) & " outputs:" & " BITSEL_u8_u1_3434_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3434_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3434_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3433_wire_constant, tmp_var);
      BITSEL_u8_u1_3434_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3444_inst flow-through 
    process(BITSEL_u8_u1_3444_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3444_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3443_wire_constant = "& Convert_SLV_To_Hex_String(konst_3443_wire_constant) & " outputs:" & " BITSEL_u8_u1_3444_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3444_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3444_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3443_wire_constant, tmp_var);
      BITSEL_u8_u1_3444_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3454_inst flow-through 
    process(BITSEL_u8_u1_3454_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3454_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3453_wire_constant = "& Convert_SLV_To_Hex_String(konst_3453_wire_constant) & " outputs:" & " BITSEL_u8_u1_3454_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3454_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3454_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3453_wire_constant, tmp_var);
      BITSEL_u8_u1_3454_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3464_inst flow-through 
    process(BITSEL_u8_u1_3464_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3464_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3463_wire_constant = "& Convert_SLV_To_Hex_String(konst_3463_wire_constant) & " outputs:" & " BITSEL_u8_u1_3464_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3464_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3464_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3463_wire_constant, tmp_var);
      BITSEL_u8_u1_3464_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3474_inst flow-through 
    process(BITSEL_u8_u1_3474_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3474_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3473_wire_constant = "& Convert_SLV_To_Hex_String(konst_3473_wire_constant) & " outputs:" & " BITSEL_u8_u1_3474_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3474_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3474_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3473_wire_constant, tmp_var);
      BITSEL_u8_u1_3474_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3484_inst flow-through 
    process(BITSEL_u8_u1_3484_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3484_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3483_wire_constant = "& Convert_SLV_To_Hex_String(konst_3483_wire_constant) & " outputs:" & " BITSEL_u8_u1_3484_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3484_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3484_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3483_wire_constant, tmp_var);
      BITSEL_u8_u1_3484_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3494_inst flow-through 
    process(BITSEL_u8_u1_3494_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3494_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3493_wire_constant = "& Convert_SLV_To_Hex_String(konst_3493_wire_constant) & " outputs:" & " BITSEL_u8_u1_3494_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3494_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3494_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3493_wire_constant, tmp_var);
      BITSEL_u8_u1_3494_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3504_inst flow-through 
    process(BITSEL_u8_u1_3504_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3504_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3503_wire_constant = "& Convert_SLV_To_Hex_String(konst_3503_wire_constant) & " outputs:" & " BITSEL_u8_u1_3504_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3504_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3504_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3503_wire_constant, tmp_var);
      BITSEL_u8_u1_3504_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3514_inst flow-through 
    process(BITSEL_u8_u1_3514_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3514_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3513_wire_constant = "& Convert_SLV_To_Hex_String(konst_3513_wire_constant) & " outputs:" & " BITSEL_u8_u1_3514_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3514_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3514_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3513_wire_constant, tmp_var);
      BITSEL_u8_u1_3514_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3524_inst flow-through 
    process(BITSEL_u8_u1_3524_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3524_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3523_wire_constant = "& Convert_SLV_To_Hex_String(konst_3523_wire_constant) & " outputs:" & " BITSEL_u8_u1_3524_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3524_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3524_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3523_wire_constant, tmp_var);
      BITSEL_u8_u1_3524_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3534_inst flow-through 
    process(BITSEL_u8_u1_3534_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3534_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3533_wire_constant = "& Convert_SLV_To_Hex_String(konst_3533_wire_constant) & " outputs:" & " BITSEL_u8_u1_3534_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3534_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3534_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3533_wire_constant, tmp_var);
      BITSEL_u8_u1_3534_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3544_inst flow-through 
    process(BITSEL_u8_u1_3544_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3544_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3543_wire_constant = "& Convert_SLV_To_Hex_String(konst_3543_wire_constant) & " outputs:" & " BITSEL_u8_u1_3544_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3544_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3544_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3543_wire_constant, tmp_var);
      BITSEL_u8_u1_3544_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3554_inst flow-through 
    process(BITSEL_u8_u1_3554_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3554_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3553_wire_constant = "& Convert_SLV_To_Hex_String(konst_3553_wire_constant) & " outputs:" & " BITSEL_u8_u1_3554_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3554_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3554_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3553_wire_constant, tmp_var);
      BITSEL_u8_u1_3554_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3564_inst flow-through 
    process(BITSEL_u8_u1_3564_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3564_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3563_wire_constant = "& Convert_SLV_To_Hex_String(konst_3563_wire_constant) & " outputs:" & " BITSEL_u8_u1_3564_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3564_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3564_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3563_wire_constant, tmp_var);
      BITSEL_u8_u1_3564_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3574_inst flow-through 
    process(BITSEL_u8_u1_3574_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3574_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3573_wire_constant = "& Convert_SLV_To_Hex_String(konst_3573_wire_constant) & " outputs:" & " BITSEL_u8_u1_3574_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3574_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3574_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3573_wire_constant, tmp_var);
      BITSEL_u8_u1_3574_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3584_inst flow-through 
    process(BITSEL_u8_u1_3584_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3584_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3583_wire_constant = "& Convert_SLV_To_Hex_String(konst_3583_wire_constant) & " outputs:" & " BITSEL_u8_u1_3584_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3584_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3584_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3583_wire_constant, tmp_var);
      BITSEL_u8_u1_3584_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3594_inst flow-through 
    process(BITSEL_u8_u1_3594_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3594_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3593_wire_constant = "& Convert_SLV_To_Hex_String(konst_3593_wire_constant) & " outputs:" & " BITSEL_u8_u1_3594_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3594_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3594_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3593_wire_constant, tmp_var);
      BITSEL_u8_u1_3594_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3602_inst flow-through 
    process(BITSEL_u8_u1_3602_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3602_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3601_wire_constant = "& Convert_SLV_To_Hex_String(konst_3601_wire_constant) & " outputs:" & " BITSEL_u8_u1_3602_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3602_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3602_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3601_wire_constant, tmp_var);
      BITSEL_u8_u1_3602_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3610_inst flow-through 
    process(BITSEL_u8_u1_3610_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3610_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3609_wire_constant = "& Convert_SLV_To_Hex_String(konst_3609_wire_constant) & " outputs:" & " BITSEL_u8_u1_3610_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3610_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3610_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3609_wire_constant, tmp_var);
      BITSEL_u8_u1_3610_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3618_inst flow-through 
    process(BITSEL_u8_u1_3618_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3618_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3617_wire_constant = "& Convert_SLV_To_Hex_String(konst_3617_wire_constant) & " outputs:" & " BITSEL_u8_u1_3618_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3618_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3618_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3617_wire_constant, tmp_var);
      BITSEL_u8_u1_3618_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3626_inst flow-through 
    process(BITSEL_u8_u1_3626_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3626_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3625_wire_constant = "& Convert_SLV_To_Hex_String(konst_3625_wire_constant) & " outputs:" & " BITSEL_u8_u1_3626_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3626_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3626_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3625_wire_constant, tmp_var);
      BITSEL_u8_u1_3626_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3634_inst flow-through 
    process(BITSEL_u8_u1_3634_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3634_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3633_wire_constant = "& Convert_SLV_To_Hex_String(konst_3633_wire_constant) & " outputs:" & " BITSEL_u8_u1_3634_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3634_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3634_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3633_wire_constant, tmp_var);
      BITSEL_u8_u1_3634_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3642_inst flow-through 
    process(BITSEL_u8_u1_3642_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3642_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3641_wire_constant = "& Convert_SLV_To_Hex_String(konst_3641_wire_constant) & " outputs:" & " BITSEL_u8_u1_3642_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3642_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3642_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3641_wire_constant, tmp_var);
      BITSEL_u8_u1_3642_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3650_inst flow-through 
    process(BITSEL_u8_u1_3650_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3650_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3649_wire_constant = "& Convert_SLV_To_Hex_String(konst_3649_wire_constant) & " outputs:" & " BITSEL_u8_u1_3650_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3650_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3650_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3649_wire_constant, tmp_var);
      BITSEL_u8_u1_3650_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3658_inst flow-through 
    process(BITSEL_u8_u1_3658_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3658_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3657_wire_constant = "& Convert_SLV_To_Hex_String(konst_3657_wire_constant) & " outputs:" & " BITSEL_u8_u1_3658_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3658_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3658_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3657_wire_constant, tmp_var);
      BITSEL_u8_u1_3658_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3666_inst flow-through 
    process(BITSEL_u8_u1_3666_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3666_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3665_wire_constant = "& Convert_SLV_To_Hex_String(konst_3665_wire_constant) & " outputs:" & " BITSEL_u8_u1_3666_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3666_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3666_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3665_wire_constant, tmp_var);
      BITSEL_u8_u1_3666_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3674_inst flow-through 
    process(BITSEL_u8_u1_3674_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3674_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3673_wire_constant = "& Convert_SLV_To_Hex_String(konst_3673_wire_constant) & " outputs:" & " BITSEL_u8_u1_3674_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3674_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3674_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3673_wire_constant, tmp_var);
      BITSEL_u8_u1_3674_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3682_inst flow-through 
    process(BITSEL_u8_u1_3682_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3682_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3681_wire_constant = "& Convert_SLV_To_Hex_String(konst_3681_wire_constant) & " outputs:" & " BITSEL_u8_u1_3682_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3682_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3682_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3681_wire_constant, tmp_var);
      BITSEL_u8_u1_3682_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3690_inst flow-through 
    process(BITSEL_u8_u1_3690_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3690_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3689_wire_constant = "& Convert_SLV_To_Hex_String(konst_3689_wire_constant) & " outputs:" & " BITSEL_u8_u1_3690_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3690_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3690_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3689_wire_constant, tmp_var);
      BITSEL_u8_u1_3690_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3698_inst flow-through 
    process(BITSEL_u8_u1_3698_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3698_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3697_wire_constant = "& Convert_SLV_To_Hex_String(konst_3697_wire_constant) & " outputs:" & " BITSEL_u8_u1_3698_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3698_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3698_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3697_wire_constant, tmp_var);
      BITSEL_u8_u1_3698_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3706_inst flow-through 
    process(BITSEL_u8_u1_3706_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3706_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3705_wire_constant = "& Convert_SLV_To_Hex_String(konst_3705_wire_constant) & " outputs:" & " BITSEL_u8_u1_3706_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3706_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3706_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3705_wire_constant, tmp_var);
      BITSEL_u8_u1_3706_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3714_inst flow-through 
    process(BITSEL_u8_u1_3714_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3714_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3713_wire_constant = "& Convert_SLV_To_Hex_String(konst_3713_wire_constant) & " outputs:" & " BITSEL_u8_u1_3714_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3714_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3714_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3713_wire_constant, tmp_var);
      BITSEL_u8_u1_3714_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3722_inst flow-through 
    process(BITSEL_u8_u1_3722_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3722_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3721_wire_constant = "& Convert_SLV_To_Hex_String(konst_3721_wire_constant) & " outputs:" & " BITSEL_u8_u1_3722_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3722_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3722_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3721_wire_constant, tmp_var);
      BITSEL_u8_u1_3722_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3730_inst flow-through 
    process(BITSEL_u8_u1_3730_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3730_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3729_wire_constant = "& Convert_SLV_To_Hex_String(konst_3729_wire_constant) & " outputs:" & " BITSEL_u8_u1_3730_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3730_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3730_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3729_wire_constant, tmp_var);
      BITSEL_u8_u1_3730_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3738_inst flow-through 
    process(BITSEL_u8_u1_3738_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3738_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3737_wire_constant = "& Convert_SLV_To_Hex_String(konst_3737_wire_constant) & " outputs:" & " BITSEL_u8_u1_3738_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3738_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3738_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3737_wire_constant, tmp_var);
      BITSEL_u8_u1_3738_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3746_inst flow-through 
    process(BITSEL_u8_u1_3746_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3746_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3745_wire_constant = "& Convert_SLV_To_Hex_String(konst_3745_wire_constant) & " outputs:" & " BITSEL_u8_u1_3746_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3746_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3746_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3745_wire_constant, tmp_var);
      BITSEL_u8_u1_3746_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3754_inst flow-through 
    process(BITSEL_u8_u1_3754_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3754_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3753_wire_constant = "& Convert_SLV_To_Hex_String(konst_3753_wire_constant) & " outputs:" & " BITSEL_u8_u1_3754_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3754_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3754_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3753_wire_constant, tmp_var);
      BITSEL_u8_u1_3754_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3762_inst flow-through 
    process(BITSEL_u8_u1_3762_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3762_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3761_wire_constant = "& Convert_SLV_To_Hex_String(konst_3761_wire_constant) & " outputs:" & " BITSEL_u8_u1_3762_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3762_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3762_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3761_wire_constant, tmp_var);
      BITSEL_u8_u1_3762_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3770_inst flow-through 
    process(BITSEL_u8_u1_3770_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3770_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3769_wire_constant = "& Convert_SLV_To_Hex_String(konst_3769_wire_constant) & " outputs:" & " BITSEL_u8_u1_3770_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3770_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3770_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3769_wire_constant, tmp_var);
      BITSEL_u8_u1_3770_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3778_inst flow-through 
    process(BITSEL_u8_u1_3778_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3778_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3777_wire_constant = "& Convert_SLV_To_Hex_String(konst_3777_wire_constant) & " outputs:" & " BITSEL_u8_u1_3778_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3778_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3778_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3777_wire_constant, tmp_var);
      BITSEL_u8_u1_3778_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3786_inst flow-through 
    process(BITSEL_u8_u1_3786_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3786_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3785_wire_constant = "& Convert_SLV_To_Hex_String(konst_3785_wire_constant) & " outputs:" & " BITSEL_u8_u1_3786_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3786_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3786_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3785_wire_constant, tmp_var);
      BITSEL_u8_u1_3786_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3794_inst flow-through 
    process(BITSEL_u8_u1_3794_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3794_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3793_wire_constant = "& Convert_SLV_To_Hex_String(konst_3793_wire_constant) & " outputs:" & " BITSEL_u8_u1_3794_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3794_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3794_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3793_wire_constant, tmp_var);
      BITSEL_u8_u1_3794_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3802_inst flow-through 
    process(BITSEL_u8_u1_3802_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3802_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3801_wire_constant = "& Convert_SLV_To_Hex_String(konst_3801_wire_constant) & " outputs:" & " BITSEL_u8_u1_3802_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3802_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3802_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3801_wire_constant, tmp_var);
      BITSEL_u8_u1_3802_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3810_inst flow-through 
    process(BITSEL_u8_u1_3810_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3810_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3809_wire_constant = "& Convert_SLV_To_Hex_String(konst_3809_wire_constant) & " outputs:" & " BITSEL_u8_u1_3810_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3810_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3810_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3809_wire_constant, tmp_var);
      BITSEL_u8_u1_3810_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3818_inst flow-through 
    process(BITSEL_u8_u1_3818_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3818_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3817_wire_constant = "& Convert_SLV_To_Hex_String(konst_3817_wire_constant) & " outputs:" & " BITSEL_u8_u1_3818_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3818_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3818_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3817_wire_constant, tmp_var);
      BITSEL_u8_u1_3818_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3826_inst flow-through 
    process(BITSEL_u8_u1_3826_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3826_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3825_wire_constant = "& Convert_SLV_To_Hex_String(konst_3825_wire_constant) & " outputs:" & " BITSEL_u8_u1_3826_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3826_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3826_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3825_wire_constant, tmp_var);
      BITSEL_u8_u1_3826_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3834_inst flow-through 
    process(BITSEL_u8_u1_3834_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3834_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3833_wire_constant = "& Convert_SLV_To_Hex_String(konst_3833_wire_constant) & " outputs:" & " BITSEL_u8_u1_3834_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3834_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3834_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3833_wire_constant, tmp_var);
      BITSEL_u8_u1_3834_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3842_inst flow-through 
    process(BITSEL_u8_u1_3842_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3842_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3841_wire_constant = "& Convert_SLV_To_Hex_String(konst_3841_wire_constant) & " outputs:" & " BITSEL_u8_u1_3842_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3842_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3842_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3841_wire_constant, tmp_var);
      BITSEL_u8_u1_3842_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3850_inst flow-through 
    process(BITSEL_u8_u1_3850_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3850_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3849_wire_constant = "& Convert_SLV_To_Hex_String(konst_3849_wire_constant) & " outputs:" & " BITSEL_u8_u1_3850_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3850_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3850_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3849_wire_constant, tmp_var);
      BITSEL_u8_u1_3850_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3858_inst flow-through 
    process(BITSEL_u8_u1_3858_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3858_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3857_wire_constant = "& Convert_SLV_To_Hex_String(konst_3857_wire_constant) & " outputs:" & " BITSEL_u8_u1_3858_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3858_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3858_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3857_wire_constant, tmp_var);
      BITSEL_u8_u1_3858_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3866_inst flow-through 
    process(BITSEL_u8_u1_3866_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3866_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3865_wire_constant = "& Convert_SLV_To_Hex_String(konst_3865_wire_constant) & " outputs:" & " BITSEL_u8_u1_3866_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3866_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3866_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3865_wire_constant, tmp_var);
      BITSEL_u8_u1_3866_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3874_inst flow-through 
    process(BITSEL_u8_u1_3874_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3874_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3873_wire_constant = "& Convert_SLV_To_Hex_String(konst_3873_wire_constant) & " outputs:" & " BITSEL_u8_u1_3874_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3874_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3874_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3873_wire_constant, tmp_var);
      BITSEL_u8_u1_3874_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3882_inst flow-through 
    process(BITSEL_u8_u1_3882_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3882_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3881_wire_constant = "& Convert_SLV_To_Hex_String(konst_3881_wire_constant) & " outputs:" & " BITSEL_u8_u1_3882_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3882_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3882_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3881_wire_constant, tmp_var);
      BITSEL_u8_u1_3882_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3890_inst flow-through 
    process(BITSEL_u8_u1_3890_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3890_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3889_wire_constant = "& Convert_SLV_To_Hex_String(konst_3889_wire_constant) & " outputs:" & " BITSEL_u8_u1_3890_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3890_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3890_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3889_wire_constant, tmp_var);
      BITSEL_u8_u1_3890_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3898_inst flow-through 
    process(BITSEL_u8_u1_3898_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3898_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3897_wire_constant = "& Convert_SLV_To_Hex_String(konst_3897_wire_constant) & " outputs:" & " BITSEL_u8_u1_3898_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3898_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3898_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3897_wire_constant, tmp_var);
      BITSEL_u8_u1_3898_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3906_inst flow-through 
    process(BITSEL_u8_u1_3906_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3906_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3905_wire_constant = "& Convert_SLV_To_Hex_String(konst_3905_wire_constant) & " outputs:" & " BITSEL_u8_u1_3906_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3906_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3906_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3905_wire_constant, tmp_var);
      BITSEL_u8_u1_3906_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3914_inst flow-through 
    process(BITSEL_u8_u1_3914_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3914_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3913_wire_constant = "& Convert_SLV_To_Hex_String(konst_3913_wire_constant) & " outputs:" & " BITSEL_u8_u1_3914_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3914_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3914_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3913_wire_constant, tmp_var);
      BITSEL_u8_u1_3914_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3922_inst flow-through 
    process(BITSEL_u8_u1_3922_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3922_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3921_wire_constant = "& Convert_SLV_To_Hex_String(konst_3921_wire_constant) & " outputs:" & " BITSEL_u8_u1_3922_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3922_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3922_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3921_wire_constant, tmp_var);
      BITSEL_u8_u1_3922_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3930_inst flow-through 
    process(BITSEL_u8_u1_3930_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3930_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3929_wire_constant = "& Convert_SLV_To_Hex_String(konst_3929_wire_constant) & " outputs:" & " BITSEL_u8_u1_3930_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3930_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3930_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3929_wire_constant, tmp_var);
      BITSEL_u8_u1_3930_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3938_inst flow-through 
    process(BITSEL_u8_u1_3938_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3938_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3937_wire_constant = "& Convert_SLV_To_Hex_String(konst_3937_wire_constant) & " outputs:" & " BITSEL_u8_u1_3938_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3938_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3938_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3937_wire_constant, tmp_var);
      BITSEL_u8_u1_3938_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3946_inst flow-through 
    process(BITSEL_u8_u1_3946_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3946_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3945_wire_constant = "& Convert_SLV_To_Hex_String(konst_3945_wire_constant) & " outputs:" & " BITSEL_u8_u1_3946_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3946_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3946_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3945_wire_constant, tmp_var);
      BITSEL_u8_u1_3946_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3954_inst flow-through 
    process(BITSEL_u8_u1_3954_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3954_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3953_wire_constant = "& Convert_SLV_To_Hex_String(konst_3953_wire_constant) & " outputs:" & " BITSEL_u8_u1_3954_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3954_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3954_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3953_wire_constant, tmp_var);
      BITSEL_u8_u1_3954_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3962_inst flow-through 
    process(BITSEL_u8_u1_3962_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3962_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3961_wire_constant = "& Convert_SLV_To_Hex_String(konst_3961_wire_constant) & " outputs:" & " BITSEL_u8_u1_3962_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3962_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3962_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3961_wire_constant, tmp_var);
      BITSEL_u8_u1_3962_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3970_inst flow-through 
    process(BITSEL_u8_u1_3970_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3970_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3969_wire_constant = "& Convert_SLV_To_Hex_String(konst_3969_wire_constant) & " outputs:" & " BITSEL_u8_u1_3970_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3970_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3970_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3969_wire_constant, tmp_var);
      BITSEL_u8_u1_3970_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3978_inst flow-through 
    process(BITSEL_u8_u1_3978_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3978_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3977_wire_constant = "& Convert_SLV_To_Hex_String(konst_3977_wire_constant) & " outputs:" & " BITSEL_u8_u1_3978_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3978_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3978_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3977_wire_constant, tmp_var);
      BITSEL_u8_u1_3978_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3986_inst flow-through 
    process(BITSEL_u8_u1_3986_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3986_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3985_wire_constant = "& Convert_SLV_To_Hex_String(konst_3985_wire_constant) & " outputs:" & " BITSEL_u8_u1_3986_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3986_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3986_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3985_wire_constant, tmp_var);
      BITSEL_u8_u1_3986_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_3994_inst flow-through 
    process(BITSEL_u8_u1_3994_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_3994_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_3993_wire_constant = "& Convert_SLV_To_Hex_String(konst_3993_wire_constant) & " outputs:" & " BITSEL_u8_u1_3994_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_3994_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_3994_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3993_wire_constant, tmp_var);
      BITSEL_u8_u1_3994_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4002_inst flow-through 
    process(BITSEL_u8_u1_4002_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_4002_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4001_wire_constant = "& Convert_SLV_To_Hex_String(konst_4001_wire_constant) & " outputs:" & " BITSEL_u8_u1_4002_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4002_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4002_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4001_wire_constant, tmp_var);
      BITSEL_u8_u1_4002_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4010_inst flow-through 
    process(BITSEL_u8_u1_4010_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_4010_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4009_wire_constant = "& Convert_SLV_To_Hex_String(konst_4009_wire_constant) & " outputs:" & " BITSEL_u8_u1_4010_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4010_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4010_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4009_wire_constant, tmp_var);
      BITSEL_u8_u1_4010_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4018_inst flow-through 
    process(BITSEL_u8_u1_4018_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_4018_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4017_wire_constant = "& Convert_SLV_To_Hex_String(konst_4017_wire_constant) & " outputs:" & " BITSEL_u8_u1_4018_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4018_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4018_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4017_wire_constant, tmp_var);
      BITSEL_u8_u1_4018_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4026_inst flow-through 
    process(BITSEL_u8_u1_4026_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_4026_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4025_wire_constant = "& Convert_SLV_To_Hex_String(konst_4025_wire_constant) & " outputs:" & " BITSEL_u8_u1_4026_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4026_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4026_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4025_wire_constant, tmp_var);
      BITSEL_u8_u1_4026_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4034_inst flow-through 
    process(BITSEL_u8_u1_4034_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_4034_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4033_wire_constant = "& Convert_SLV_To_Hex_String(konst_4033_wire_constant) & " outputs:" & " BITSEL_u8_u1_4034_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4034_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4034_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4033_wire_constant, tmp_var);
      BITSEL_u8_u1_4034_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4042_inst flow-through 
    process(BITSEL_u8_u1_4042_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_4042_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4041_wire_constant = "& Convert_SLV_To_Hex_String(konst_4041_wire_constant) & " outputs:" & " BITSEL_u8_u1_4042_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4042_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4042_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4041_wire_constant, tmp_var);
      BITSEL_u8_u1_4042_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4050_inst flow-through 
    process(BITSEL_u8_u1_4050_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_4050_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4049_wire_constant = "& Convert_SLV_To_Hex_String(konst_4049_wire_constant) & " outputs:" & " BITSEL_u8_u1_4050_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4050_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4050_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4049_wire_constant, tmp_var);
      BITSEL_u8_u1_4050_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4058_inst flow-through 
    process(BITSEL_u8_u1_4058_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_4058_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4057_wire_constant = "& Convert_SLV_To_Hex_String(konst_4057_wire_constant) & " outputs:" & " BITSEL_u8_u1_4058_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4058_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4058_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4057_wire_constant, tmp_var);
      BITSEL_u8_u1_4058_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4066_inst flow-through 
    process(BITSEL_u8_u1_4066_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_4066_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4065_wire_constant = "& Convert_SLV_To_Hex_String(konst_4065_wire_constant) & " outputs:" & " BITSEL_u8_u1_4066_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4066_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4066_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4065_wire_constant, tmp_var);
      BITSEL_u8_u1_4066_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4074_inst flow-through 
    process(BITSEL_u8_u1_4074_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_4074_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4073_wire_constant = "& Convert_SLV_To_Hex_String(konst_4073_wire_constant) & " outputs:" & " BITSEL_u8_u1_4074_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4074_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4074_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4073_wire_constant, tmp_var);
      BITSEL_u8_u1_4074_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4082_inst flow-through 
    process(BITSEL_u8_u1_4082_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_4082_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4081_wire_constant = "& Convert_SLV_To_Hex_String(konst_4081_wire_constant) & " outputs:" & " BITSEL_u8_u1_4082_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4082_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4082_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4081_wire_constant, tmp_var);
      BITSEL_u8_u1_4082_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4090_inst flow-through 
    process(BITSEL_u8_u1_4090_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_4090_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4089_wire_constant = "& Convert_SLV_To_Hex_String(konst_4089_wire_constant) & " outputs:" & " BITSEL_u8_u1_4090_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4090_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4090_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4089_wire_constant, tmp_var);
      BITSEL_u8_u1_4090_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4098_inst flow-through 
    process(BITSEL_u8_u1_4098_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_4098_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4097_wire_constant = "& Convert_SLV_To_Hex_String(konst_4097_wire_constant) & " outputs:" & " BITSEL_u8_u1_4098_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4098_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4098_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4097_wire_constant, tmp_var);
      BITSEL_u8_u1_4098_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4106_inst flow-through 
    process(BITSEL_u8_u1_4106_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_4106_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4105_wire_constant = "& Convert_SLV_To_Hex_String(konst_4105_wire_constant) & " outputs:" & " BITSEL_u8_u1_4106_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4106_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4106_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4105_wire_constant, tmp_var);
      BITSEL_u8_u1_4106_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4114_inst flow-through 
    process(BITSEL_u8_u1_4114_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_4114_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4113_wire_constant = "& Convert_SLV_To_Hex_String(konst_4113_wire_constant) & " outputs:" & " BITSEL_u8_u1_4114_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4114_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4114_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4113_wire_constant, tmp_var);
      BITSEL_u8_u1_4114_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4122_inst flow-through 
    process(BITSEL_u8_u1_4122_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_4122_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4121_wire_constant = "& Convert_SLV_To_Hex_String(konst_4121_wire_constant) & " outputs:" & " BITSEL_u8_u1_4122_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4122_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4122_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4121_wire_constant, tmp_var);
      BITSEL_u8_u1_4122_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4130_inst flow-through 
    process(BITSEL_u8_u1_4130_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_4130_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4129_wire_constant = "& Convert_SLV_To_Hex_String(konst_4129_wire_constant) & " outputs:" & " BITSEL_u8_u1_4130_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4130_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4130_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4129_wire_constant, tmp_var);
      BITSEL_u8_u1_4130_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4138_inst flow-through 
    process(BITSEL_u8_u1_4138_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_4138_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4137_wire_constant = "& Convert_SLV_To_Hex_String(konst_4137_wire_constant) & " outputs:" & " BITSEL_u8_u1_4138_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4138_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4138_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4137_wire_constant, tmp_var);
      BITSEL_u8_u1_4138_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4146_inst flow-through 
    process(BITSEL_u8_u1_4146_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_4146_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4145_wire_constant = "& Convert_SLV_To_Hex_String(konst_4145_wire_constant) & " outputs:" & " BITSEL_u8_u1_4146_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4146_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4146_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4145_wire_constant, tmp_var);
      BITSEL_u8_u1_4146_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4154_inst flow-through 
    process(BITSEL_u8_u1_4154_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_4154_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4153_wire_constant = "& Convert_SLV_To_Hex_String(konst_4153_wire_constant) & " outputs:" & " BITSEL_u8_u1_4154_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4154_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4154_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4153_wire_constant, tmp_var);
      BITSEL_u8_u1_4154_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4162_inst flow-through 
    process(BITSEL_u8_u1_4162_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_4162_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4161_wire_constant = "& Convert_SLV_To_Hex_String(konst_4161_wire_constant) & " outputs:" & " BITSEL_u8_u1_4162_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4162_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4162_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4161_wire_constant, tmp_var);
      BITSEL_u8_u1_4162_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4170_inst flow-through 
    process(BITSEL_u8_u1_4170_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_4170_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4169_wire_constant = "& Convert_SLV_To_Hex_String(konst_4169_wire_constant) & " outputs:" & " BITSEL_u8_u1_4170_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4170_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4170_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4169_wire_constant, tmp_var);
      BITSEL_u8_u1_4170_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4178_inst flow-through 
    process(BITSEL_u8_u1_4178_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_4178_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4177_wire_constant = "& Convert_SLV_To_Hex_String(konst_4177_wire_constant) & " outputs:" & " BITSEL_u8_u1_4178_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4178_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4178_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4177_wire_constant, tmp_var);
      BITSEL_u8_u1_4178_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4186_inst flow-through 
    process(BITSEL_u8_u1_4186_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_4186_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4185_wire_constant = "& Convert_SLV_To_Hex_String(konst_4185_wire_constant) & " outputs:" & " BITSEL_u8_u1_4186_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4186_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4186_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4185_wire_constant, tmp_var);
      BITSEL_u8_u1_4186_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4194_inst flow-through 
    process(BITSEL_u8_u1_4194_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_4194_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4193_wire_constant = "& Convert_SLV_To_Hex_String(konst_4193_wire_constant) & " outputs:" & " BITSEL_u8_u1_4194_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4194_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4194_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4193_wire_constant, tmp_var);
      BITSEL_u8_u1_4194_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4202_inst flow-through 
    process(BITSEL_u8_u1_4202_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_4202_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4201_wire_constant = "& Convert_SLV_To_Hex_String(konst_4201_wire_constant) & " outputs:" & " BITSEL_u8_u1_4202_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4202_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4202_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4201_wire_constant, tmp_var);
      BITSEL_u8_u1_4202_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4210_inst flow-through 
    process(BITSEL_u8_u1_4210_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_4210_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4209_wire_constant = "& Convert_SLV_To_Hex_String(konst_4209_wire_constant) & " outputs:" & " BITSEL_u8_u1_4210_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4210_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4210_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4209_wire_constant, tmp_var);
      BITSEL_u8_u1_4210_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4218_inst flow-through 
    process(BITSEL_u8_u1_4218_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_4218_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4217_wire_constant = "& Convert_SLV_To_Hex_String(konst_4217_wire_constant) & " outputs:" & " BITSEL_u8_u1_4218_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4218_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4218_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4217_wire_constant, tmp_var);
      BITSEL_u8_u1_4218_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4226_inst flow-through 
    process(BITSEL_u8_u1_4226_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_4226_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4225_wire_constant = "& Convert_SLV_To_Hex_String(konst_4225_wire_constant) & " outputs:" & " BITSEL_u8_u1_4226_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4226_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4226_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4225_wire_constant, tmp_var);
      BITSEL_u8_u1_4226_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4234_inst flow-through 
    process(BITSEL_u8_u1_4234_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_4234_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4233_wire_constant = "& Convert_SLV_To_Hex_String(konst_4233_wire_constant) & " outputs:" & " BITSEL_u8_u1_4234_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4234_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4234_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4233_wire_constant, tmp_var);
      BITSEL_u8_u1_4234_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4242_inst flow-through 
    process(BITSEL_u8_u1_4242_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_4242_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4241_wire_constant = "& Convert_SLV_To_Hex_String(konst_4241_wire_constant) & " outputs:" & " BITSEL_u8_u1_4242_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4242_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4242_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4241_wire_constant, tmp_var);
      BITSEL_u8_u1_4242_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4250_inst flow-through 
    process(BITSEL_u8_u1_4250_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_4250_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4249_wire_constant = "& Convert_SLV_To_Hex_String(konst_4249_wire_constant) & " outputs:" & " BITSEL_u8_u1_4250_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4250_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4250_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4249_wire_constant, tmp_var);
      BITSEL_u8_u1_4250_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4258_inst flow-through 
    process(BITSEL_u8_u1_4258_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_4258_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4257_wire_constant = "& Convert_SLV_To_Hex_String(konst_4257_wire_constant) & " outputs:" & " BITSEL_u8_u1_4258_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4258_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4258_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4257_wire_constant, tmp_var);
      BITSEL_u8_u1_4258_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4266_inst flow-through 
    process(BITSEL_u8_u1_4266_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_4266_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4265_wire_constant = "& Convert_SLV_To_Hex_String(konst_4265_wire_constant) & " outputs:" & " BITSEL_u8_u1_4266_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4266_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4266_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4265_wire_constant, tmp_var);
      BITSEL_u8_u1_4266_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4274_inst flow-through 
    process(BITSEL_u8_u1_4274_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_4274_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4273_wire_constant = "& Convert_SLV_To_Hex_String(konst_4273_wire_constant) & " outputs:" & " BITSEL_u8_u1_4274_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4274_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4274_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4273_wire_constant, tmp_var);
      BITSEL_u8_u1_4274_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4282_inst flow-through 
    process(BITSEL_u8_u1_4282_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_4282_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4281_wire_constant = "& Convert_SLV_To_Hex_String(konst_4281_wire_constant) & " outputs:" & " BITSEL_u8_u1_4282_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4282_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4282_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4281_wire_constant, tmp_var);
      BITSEL_u8_u1_4282_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4290_inst flow-through 
    process(BITSEL_u8_u1_4290_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_4290_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4289_wire_constant = "& Convert_SLV_To_Hex_String(konst_4289_wire_constant) & " outputs:" & " BITSEL_u8_u1_4290_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4290_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4290_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4289_wire_constant, tmp_var);
      BITSEL_u8_u1_4290_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4298_inst flow-through 
    process(BITSEL_u8_u1_4298_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_4298_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4297_wire_constant = "& Convert_SLV_To_Hex_String(konst_4297_wire_constant) & " outputs:" & " BITSEL_u8_u1_4298_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4298_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4298_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4297_wire_constant, tmp_var);
      BITSEL_u8_u1_4298_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4306_inst flow-through 
    process(BITSEL_u8_u1_4306_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_4306_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4305_wire_constant = "& Convert_SLV_To_Hex_String(konst_4305_wire_constant) & " outputs:" & " BITSEL_u8_u1_4306_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4306_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4306_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4305_wire_constant, tmp_var);
      BITSEL_u8_u1_4306_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4314_inst flow-through 
    process(BITSEL_u8_u1_4314_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_4314_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4313_wire_constant = "& Convert_SLV_To_Hex_String(konst_4313_wire_constant) & " outputs:" & " BITSEL_u8_u1_4314_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4314_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4314_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4313_wire_constant, tmp_var);
      BITSEL_u8_u1_4314_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4322_inst flow-through 
    process(BITSEL_u8_u1_4322_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_4322_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4321_wire_constant = "& Convert_SLV_To_Hex_String(konst_4321_wire_constant) & " outputs:" & " BITSEL_u8_u1_4322_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4322_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4322_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4321_wire_constant, tmp_var);
      BITSEL_u8_u1_4322_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4330_inst flow-through 
    process(BITSEL_u8_u1_4330_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_4330_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4329_wire_constant = "& Convert_SLV_To_Hex_String(konst_4329_wire_constant) & " outputs:" & " BITSEL_u8_u1_4330_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4330_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4330_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4329_wire_constant, tmp_var);
      BITSEL_u8_u1_4330_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4338_inst flow-through 
    process(BITSEL_u8_u1_4338_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_4338_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4337_wire_constant = "& Convert_SLV_To_Hex_String(konst_4337_wire_constant) & " outputs:" & " BITSEL_u8_u1_4338_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4338_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4338_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4337_wire_constant, tmp_var);
      BITSEL_u8_u1_4338_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4346_inst flow-through 
    process(BITSEL_u8_u1_4346_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_4346_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4345_wire_constant = "& Convert_SLV_To_Hex_String(konst_4345_wire_constant) & " outputs:" & " BITSEL_u8_u1_4346_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4346_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4346_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4345_wire_constant, tmp_var);
      BITSEL_u8_u1_4346_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4354_inst flow-through 
    process(BITSEL_u8_u1_4354_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_4354_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4353_wire_constant = "& Convert_SLV_To_Hex_String(konst_4353_wire_constant) & " outputs:" & " BITSEL_u8_u1_4354_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4354_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4354_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4353_wire_constant, tmp_var);
      BITSEL_u8_u1_4354_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4362_inst flow-through 
    process(BITSEL_u8_u1_4362_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_4362_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4361_wire_constant = "& Convert_SLV_To_Hex_String(konst_4361_wire_constant) & " outputs:" & " BITSEL_u8_u1_4362_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4362_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4362_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4361_wire_constant, tmp_var);
      BITSEL_u8_u1_4362_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4370_inst flow-through 
    process(BITSEL_u8_u1_4370_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_4370_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4369_wire_constant = "& Convert_SLV_To_Hex_String(konst_4369_wire_constant) & " outputs:" & " BITSEL_u8_u1_4370_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4370_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4370_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4369_wire_constant, tmp_var);
      BITSEL_u8_u1_4370_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4378_inst flow-through 
    process(BITSEL_u8_u1_4378_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_4378_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4377_wire_constant = "& Convert_SLV_To_Hex_String(konst_4377_wire_constant) & " outputs:" & " BITSEL_u8_u1_4378_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4378_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4378_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4377_wire_constant, tmp_var);
      BITSEL_u8_u1_4378_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4386_inst flow-through 
    process(BITSEL_u8_u1_4386_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_4386_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4385_wire_constant = "& Convert_SLV_To_Hex_String(konst_4385_wire_constant) & " outputs:" & " BITSEL_u8_u1_4386_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4386_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4386_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4385_wire_constant, tmp_var);
      BITSEL_u8_u1_4386_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4394_inst flow-through 
    process(BITSEL_u8_u1_4394_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_4394_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4393_wire_constant = "& Convert_SLV_To_Hex_String(konst_4393_wire_constant) & " outputs:" & " BITSEL_u8_u1_4394_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4394_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4394_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4393_wire_constant, tmp_var);
      BITSEL_u8_u1_4394_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4402_inst flow-through 
    process(BITSEL_u8_u1_4402_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_4402_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4401_wire_constant = "& Convert_SLV_To_Hex_String(konst_4401_wire_constant) & " outputs:" & " BITSEL_u8_u1_4402_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4402_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4402_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4401_wire_constant, tmp_var);
      BITSEL_u8_u1_4402_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4410_inst flow-through 
    process(BITSEL_u8_u1_4410_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_4410_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4409_wire_constant = "& Convert_SLV_To_Hex_String(konst_4409_wire_constant) & " outputs:" & " BITSEL_u8_u1_4410_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4410_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4410_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4409_wire_constant, tmp_var);
      BITSEL_u8_u1_4410_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4418_inst flow-through 
    process(BITSEL_u8_u1_4418_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_4418_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4417_wire_constant = "& Convert_SLV_To_Hex_String(konst_4417_wire_constant) & " outputs:" & " BITSEL_u8_u1_4418_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4418_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4418_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4417_wire_constant, tmp_var);
      BITSEL_u8_u1_4418_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4426_inst flow-through 
    process(BITSEL_u8_u1_4426_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_4426_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4425_wire_constant = "& Convert_SLV_To_Hex_String(konst_4425_wire_constant) & " outputs:" & " BITSEL_u8_u1_4426_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4426_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4426_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4425_wire_constant, tmp_var);
      BITSEL_u8_u1_4426_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4434_inst flow-through 
    process(BITSEL_u8_u1_4434_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_4434_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4433_wire_constant = "& Convert_SLV_To_Hex_String(konst_4433_wire_constant) & " outputs:" & " BITSEL_u8_u1_4434_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4434_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4434_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4433_wire_constant, tmp_var);
      BITSEL_u8_u1_4434_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4442_inst flow-through 
    process(BITSEL_u8_u1_4442_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_4442_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4441_wire_constant = "& Convert_SLV_To_Hex_String(konst_4441_wire_constant) & " outputs:" & " BITSEL_u8_u1_4442_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4442_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4442_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4441_wire_constant, tmp_var);
      BITSEL_u8_u1_4442_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4450_inst flow-through 
    process(BITSEL_u8_u1_4450_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_4450_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4449_wire_constant = "& Convert_SLV_To_Hex_String(konst_4449_wire_constant) & " outputs:" & " BITSEL_u8_u1_4450_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4450_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4450_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4449_wire_constant, tmp_var);
      BITSEL_u8_u1_4450_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4458_inst flow-through 
    process(BITSEL_u8_u1_4458_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_4458_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4457_wire_constant = "& Convert_SLV_To_Hex_String(konst_4457_wire_constant) & " outputs:" & " BITSEL_u8_u1_4458_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4458_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4458_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4457_wire_constant, tmp_var);
      BITSEL_u8_u1_4458_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4466_inst flow-through 
    process(BITSEL_u8_u1_4466_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_4466_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4465_wire_constant = "& Convert_SLV_To_Hex_String(konst_4465_wire_constant) & " outputs:" & " BITSEL_u8_u1_4466_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4466_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4466_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4465_wire_constant, tmp_var);
      BITSEL_u8_u1_4466_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4474_inst flow-through 
    process(BITSEL_u8_u1_4474_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_4474_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4473_wire_constant = "& Convert_SLV_To_Hex_String(konst_4473_wire_constant) & " outputs:" & " BITSEL_u8_u1_4474_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4474_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4474_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4473_wire_constant, tmp_var);
      BITSEL_u8_u1_4474_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4482_inst flow-through 
    process(BITSEL_u8_u1_4482_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_4482_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4481_wire_constant = "& Convert_SLV_To_Hex_String(konst_4481_wire_constant) & " outputs:" & " BITSEL_u8_u1_4482_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4482_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4482_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4481_wire_constant, tmp_var);
      BITSEL_u8_u1_4482_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4490_inst flow-through 
    process(BITSEL_u8_u1_4490_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_4490_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4489_wire_constant = "& Convert_SLV_To_Hex_String(konst_4489_wire_constant) & " outputs:" & " BITSEL_u8_u1_4490_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4490_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4490_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4489_wire_constant, tmp_var);
      BITSEL_u8_u1_4490_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4498_inst flow-through 
    process(BITSEL_u8_u1_4498_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_4498_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4497_wire_constant = "& Convert_SLV_To_Hex_String(konst_4497_wire_constant) & " outputs:" & " BITSEL_u8_u1_4498_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4498_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4498_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4497_wire_constant, tmp_var);
      BITSEL_u8_u1_4498_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4506_inst flow-through 
    process(BITSEL_u8_u1_4506_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_4506_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4505_wire_constant = "& Convert_SLV_To_Hex_String(konst_4505_wire_constant) & " outputs:" & " BITSEL_u8_u1_4506_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4506_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4506_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4505_wire_constant, tmp_var);
      BITSEL_u8_u1_4506_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4514_inst flow-through 
    process(BITSEL_u8_u1_4514_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_4514_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4513_wire_constant = "& Convert_SLV_To_Hex_String(konst_4513_wire_constant) & " outputs:" & " BITSEL_u8_u1_4514_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4514_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4514_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4513_wire_constant, tmp_var);
      BITSEL_u8_u1_4514_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4522_inst flow-through 
    process(BITSEL_u8_u1_4522_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_4522_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4521_wire_constant = "& Convert_SLV_To_Hex_String(konst_4521_wire_constant) & " outputs:" & " BITSEL_u8_u1_4522_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4522_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4522_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4521_wire_constant, tmp_var);
      BITSEL_u8_u1_4522_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4530_inst flow-through 
    process(BITSEL_u8_u1_4530_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_4530_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4529_wire_constant = "& Convert_SLV_To_Hex_String(konst_4529_wire_constant) & " outputs:" & " BITSEL_u8_u1_4530_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4530_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4530_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4529_wire_constant, tmp_var);
      BITSEL_u8_u1_4530_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4538_inst flow-through 
    process(BITSEL_u8_u1_4538_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_4538_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4537_wire_constant = "& Convert_SLV_To_Hex_String(konst_4537_wire_constant) & " outputs:" & " BITSEL_u8_u1_4538_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4538_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4538_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4537_wire_constant, tmp_var);
      BITSEL_u8_u1_4538_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4546_inst flow-through 
    process(BITSEL_u8_u1_4546_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_4546_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4545_wire_constant = "& Convert_SLV_To_Hex_String(konst_4545_wire_constant) & " outputs:" & " BITSEL_u8_u1_4546_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4546_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4546_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4545_wire_constant, tmp_var);
      BITSEL_u8_u1_4546_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4554_inst flow-through 
    process(BITSEL_u8_u1_4554_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_4554_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4553_wire_constant = "& Convert_SLV_To_Hex_String(konst_4553_wire_constant) & " outputs:" & " BITSEL_u8_u1_4554_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4554_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4554_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4553_wire_constant, tmp_var);
      BITSEL_u8_u1_4554_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4562_inst flow-through 
    process(BITSEL_u8_u1_4562_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_4562_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4561_wire_constant = "& Convert_SLV_To_Hex_String(konst_4561_wire_constant) & " outputs:" & " BITSEL_u8_u1_4562_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4562_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4562_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4561_wire_constant, tmp_var);
      BITSEL_u8_u1_4562_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4570_inst flow-through 
    process(BITSEL_u8_u1_4570_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_4570_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4569_wire_constant = "& Convert_SLV_To_Hex_String(konst_4569_wire_constant) & " outputs:" & " BITSEL_u8_u1_4570_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4570_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4570_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4569_wire_constant, tmp_var);
      BITSEL_u8_u1_4570_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4578_inst flow-through 
    process(BITSEL_u8_u1_4578_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_4578_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4577_wire_constant = "& Convert_SLV_To_Hex_String(konst_4577_wire_constant) & " outputs:" & " BITSEL_u8_u1_4578_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4578_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4578_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4577_wire_constant, tmp_var);
      BITSEL_u8_u1_4578_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4586_inst flow-through 
    process(BITSEL_u8_u1_4586_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_4586_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4585_wire_constant = "& Convert_SLV_To_Hex_String(konst_4585_wire_constant) & " outputs:" & " BITSEL_u8_u1_4586_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4586_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4586_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4585_wire_constant, tmp_var);
      BITSEL_u8_u1_4586_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4594_inst flow-through 
    process(BITSEL_u8_u1_4594_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_4594_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4593_wire_constant = "& Convert_SLV_To_Hex_String(konst_4593_wire_constant) & " outputs:" & " BITSEL_u8_u1_4594_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4594_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4594_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4593_wire_constant, tmp_var);
      BITSEL_u8_u1_4594_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4602_inst flow-through 
    process(BITSEL_u8_u1_4602_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_2:DP:BITSEL_u8_u1_4602_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4601_wire_constant = "& Convert_SLV_To_Hex_String(konst_4601_wire_constant) & " outputs:" & " BITSEL_u8_u1_4602_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4602_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4602_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4601_wire_constant, tmp_var);
      BITSEL_u8_u1_4602_wire <= tmp_var; -- 
    end process;
    -- 
  end Block; -- data_path
  -- 
end Inv_Sbox_2_Volatile_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library GhdlLink;
use GhdlLink.LogUtilities.all;
library work;
use work.ahir_system_global_package.all;
entity Inv_Sbox_3_Volatile is -- 
  port ( -- 
    clk, reset: in std_logic; 
    s_in : in  std_logic_vector(7 downto 0);
    s_out : out  std_logic_vector(7 downto 0)-- 
  );
  -- 
end entity Inv_Sbox_3_Volatile;
architecture Inv_Sbox_3_Volatile_arch of Inv_Sbox_3_Volatile is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector(8-1 downto 0);
  signal default_zero_sig: std_logic;
  -- input port buffer signals
  signal s_in_buffer :  std_logic_vector(7 downto 0);
  -- output port buffer signals
  signal s_out_buffer :  std_logic_vector(7 downto 0);
  -- volatile/operator module components. 
  signal global_clock_cycle_count: integer := 0;
  -- 
begin --  
  ---------------------------------------------------------- 
  process(clk)  
  begin -- 
    if(clk'event and clk = '1') then -- 
      if(reset = '1') then -- 
        global_clock_cycle_count <= 0; --
      else -- 
        global_clock_cycle_count <= global_clock_cycle_count + 1; -- 
      end if; --
    end if; --
  end process;
  ---------------------------------------------------------- 
  -- input handling ------------------------------------------------
  s_in_buffer <= s_in;
  -- output handling  -------------------------------------------------------
  s_out <= s_out_buffer;
  -- the control path --------------------------------------------------
  default_zero_sig <= '0';
  -- volatile module, no control path
  -- the data path
  data_path: Block -- 
    signal BITSEL_u8_u1_4614_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4624_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4634_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4644_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4654_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4664_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4674_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4684_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4694_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4704_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4714_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4724_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4734_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4744_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4754_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4764_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4774_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4784_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4794_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4804_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4814_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4824_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4834_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4844_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4854_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4864_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4874_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4884_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4894_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4904_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4914_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4924_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4934_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4944_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4954_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4964_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4974_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4984_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4994_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5004_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5014_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5024_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5034_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5044_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5054_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5064_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5074_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5084_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5094_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5104_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5114_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5124_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5134_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5144_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5154_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5164_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5174_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5184_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5194_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5204_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5214_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5224_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5234_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5244_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5254_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5264_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5274_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5284_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5294_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5304_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5314_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5324_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5334_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5344_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5354_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5364_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5374_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5384_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5394_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5404_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5414_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5424_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5434_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5444_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5454_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5464_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5474_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5484_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5494_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5504_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5514_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5524_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5534_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5544_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5554_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5564_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5574_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5584_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5594_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5604_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5614_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5624_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5634_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5644_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5654_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5664_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5674_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5684_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5694_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5704_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5714_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5724_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5734_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5744_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5754_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5764_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5774_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5784_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5794_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5804_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5814_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5824_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5834_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5844_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5854_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5864_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5874_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5884_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5894_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5902_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5910_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5918_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5926_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5934_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5942_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5950_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5958_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5966_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5974_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5982_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5990_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5998_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6006_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6014_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6022_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6030_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6038_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6046_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6054_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6062_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6070_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6078_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6086_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6094_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6102_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6110_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6118_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6126_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6134_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6142_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6150_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6158_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6166_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6174_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6182_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6190_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6198_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6206_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6214_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6222_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6230_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6238_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6246_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6254_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6262_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6270_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6278_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6286_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6294_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6302_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6310_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6318_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6326_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6334_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6342_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6350_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6358_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6366_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6374_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6382_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6390_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6398_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6406_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6414_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6422_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6430_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6438_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6446_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6454_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6462_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6470_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6478_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6486_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6494_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6502_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6510_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6518_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6526_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6534_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6542_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6550_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6558_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6566_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6574_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6582_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6590_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6598_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6606_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6614_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6622_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6630_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6638_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6646_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6654_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6662_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6670_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6678_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6686_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6694_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6702_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6710_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6718_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6726_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6734_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6742_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6750_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6758_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6766_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6774_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6782_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6790_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6798_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6806_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6814_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6822_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6830_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6838_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6846_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6854_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6862_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6870_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6878_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6886_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6894_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6902_wire : std_logic_vector(0 downto 0);
    signal IMA0_4620 : std_logic_vector(7 downto 0);
    signal IMA100_5620 : std_logic_vector(7 downto 0);
    signal IMA101_5630 : std_logic_vector(7 downto 0);
    signal IMA102_5640 : std_logic_vector(7 downto 0);
    signal IMA103_5650 : std_logic_vector(7 downto 0);
    signal IMA104_5660 : std_logic_vector(7 downto 0);
    signal IMA105_5670 : std_logic_vector(7 downto 0);
    signal IMA106_5680 : std_logic_vector(7 downto 0);
    signal IMA107_5690 : std_logic_vector(7 downto 0);
    signal IMA108_5700 : std_logic_vector(7 downto 0);
    signal IMA109_5710 : std_logic_vector(7 downto 0);
    signal IMA10_4720 : std_logic_vector(7 downto 0);
    signal IMA110_5720 : std_logic_vector(7 downto 0);
    signal IMA111_5730 : std_logic_vector(7 downto 0);
    signal IMA112_5740 : std_logic_vector(7 downto 0);
    signal IMA113_5750 : std_logic_vector(7 downto 0);
    signal IMA114_5760 : std_logic_vector(7 downto 0);
    signal IMA115_5770 : std_logic_vector(7 downto 0);
    signal IMA116_5780 : std_logic_vector(7 downto 0);
    signal IMA117_5790 : std_logic_vector(7 downto 0);
    signal IMA118_5800 : std_logic_vector(7 downto 0);
    signal IMA119_5810 : std_logic_vector(7 downto 0);
    signal IMA11_4730 : std_logic_vector(7 downto 0);
    signal IMA120_5820 : std_logic_vector(7 downto 0);
    signal IMA121_5830 : std_logic_vector(7 downto 0);
    signal IMA122_5840 : std_logic_vector(7 downto 0);
    signal IMA123_5850 : std_logic_vector(7 downto 0);
    signal IMA124_5860 : std_logic_vector(7 downto 0);
    signal IMA125_5870 : std_logic_vector(7 downto 0);
    signal IMA126_5880 : std_logic_vector(7 downto 0);
    signal IMA127_5890 : std_logic_vector(7 downto 0);
    signal IMA12_4740 : std_logic_vector(7 downto 0);
    signal IMA13_4750 : std_logic_vector(7 downto 0);
    signal IMA14_4760 : std_logic_vector(7 downto 0);
    signal IMA15_4770 : std_logic_vector(7 downto 0);
    signal IMA16_4780 : std_logic_vector(7 downto 0);
    signal IMA17_4790 : std_logic_vector(7 downto 0);
    signal IMA18_4800 : std_logic_vector(7 downto 0);
    signal IMA19_4810 : std_logic_vector(7 downto 0);
    signal IMA1_4630 : std_logic_vector(7 downto 0);
    signal IMA20_4820 : std_logic_vector(7 downto 0);
    signal IMA21_4830 : std_logic_vector(7 downto 0);
    signal IMA22_4840 : std_logic_vector(7 downto 0);
    signal IMA23_4850 : std_logic_vector(7 downto 0);
    signal IMA24_4860 : std_logic_vector(7 downto 0);
    signal IMA25_4870 : std_logic_vector(7 downto 0);
    signal IMA26_4880 : std_logic_vector(7 downto 0);
    signal IMA27_4890 : std_logic_vector(7 downto 0);
    signal IMA28_4900 : std_logic_vector(7 downto 0);
    signal IMA29_4910 : std_logic_vector(7 downto 0);
    signal IMA2_4640 : std_logic_vector(7 downto 0);
    signal IMA30_4920 : std_logic_vector(7 downto 0);
    signal IMA31_4930 : std_logic_vector(7 downto 0);
    signal IMA32_4940 : std_logic_vector(7 downto 0);
    signal IMA33_4950 : std_logic_vector(7 downto 0);
    signal IMA34_4960 : std_logic_vector(7 downto 0);
    signal IMA35_4970 : std_logic_vector(7 downto 0);
    signal IMA36_4980 : std_logic_vector(7 downto 0);
    signal IMA37_4990 : std_logic_vector(7 downto 0);
    signal IMA38_5000 : std_logic_vector(7 downto 0);
    signal IMA39_5010 : std_logic_vector(7 downto 0);
    signal IMA3_4650 : std_logic_vector(7 downto 0);
    signal IMA40_5020 : std_logic_vector(7 downto 0);
    signal IMA41_5030 : std_logic_vector(7 downto 0);
    signal IMA42_5040 : std_logic_vector(7 downto 0);
    signal IMA43_5050 : std_logic_vector(7 downto 0);
    signal IMA44_5060 : std_logic_vector(7 downto 0);
    signal IMA45_5070 : std_logic_vector(7 downto 0);
    signal IMA46_5080 : std_logic_vector(7 downto 0);
    signal IMA47_5090 : std_logic_vector(7 downto 0);
    signal IMA48_5100 : std_logic_vector(7 downto 0);
    signal IMA49_5110 : std_logic_vector(7 downto 0);
    signal IMA4_4660 : std_logic_vector(7 downto 0);
    signal IMA50_5120 : std_logic_vector(7 downto 0);
    signal IMA51_5130 : std_logic_vector(7 downto 0);
    signal IMA52_5140 : std_logic_vector(7 downto 0);
    signal IMA53_5150 : std_logic_vector(7 downto 0);
    signal IMA54_5160 : std_logic_vector(7 downto 0);
    signal IMA55_5170 : std_logic_vector(7 downto 0);
    signal IMA56_5180 : std_logic_vector(7 downto 0);
    signal IMA57_5190 : std_logic_vector(7 downto 0);
    signal IMA58_5200 : std_logic_vector(7 downto 0);
    signal IMA59_5210 : std_logic_vector(7 downto 0);
    signal IMA5_4670 : std_logic_vector(7 downto 0);
    signal IMA60_5220 : std_logic_vector(7 downto 0);
    signal IMA61_5230 : std_logic_vector(7 downto 0);
    signal IMA62_5240 : std_logic_vector(7 downto 0);
    signal IMA63_5250 : std_logic_vector(7 downto 0);
    signal IMA64_5260 : std_logic_vector(7 downto 0);
    signal IMA65_5270 : std_logic_vector(7 downto 0);
    signal IMA66_5280 : std_logic_vector(7 downto 0);
    signal IMA67_5290 : std_logic_vector(7 downto 0);
    signal IMA68_5300 : std_logic_vector(7 downto 0);
    signal IMA69_5310 : std_logic_vector(7 downto 0);
    signal IMA6_4680 : std_logic_vector(7 downto 0);
    signal IMA70_5320 : std_logic_vector(7 downto 0);
    signal IMA71_5330 : std_logic_vector(7 downto 0);
    signal IMA72_5340 : std_logic_vector(7 downto 0);
    signal IMA73_5350 : std_logic_vector(7 downto 0);
    signal IMA74_5360 : std_logic_vector(7 downto 0);
    signal IMA75_5370 : std_logic_vector(7 downto 0);
    signal IMA76_5380 : std_logic_vector(7 downto 0);
    signal IMA77_5390 : std_logic_vector(7 downto 0);
    signal IMA78_5400 : std_logic_vector(7 downto 0);
    signal IMA79_5410 : std_logic_vector(7 downto 0);
    signal IMA7_4690 : std_logic_vector(7 downto 0);
    signal IMA80_5420 : std_logic_vector(7 downto 0);
    signal IMA81_5430 : std_logic_vector(7 downto 0);
    signal IMA82_5440 : std_logic_vector(7 downto 0);
    signal IMA83_5450 : std_logic_vector(7 downto 0);
    signal IMA84_5460 : std_logic_vector(7 downto 0);
    signal IMA85_5470 : std_logic_vector(7 downto 0);
    signal IMA86_5480 : std_logic_vector(7 downto 0);
    signal IMA87_5490 : std_logic_vector(7 downto 0);
    signal IMA88_5500 : std_logic_vector(7 downto 0);
    signal IMA89_5510 : std_logic_vector(7 downto 0);
    signal IMA8_4700 : std_logic_vector(7 downto 0);
    signal IMA90_5520 : std_logic_vector(7 downto 0);
    signal IMA91_5530 : std_logic_vector(7 downto 0);
    signal IMA92_5540 : std_logic_vector(7 downto 0);
    signal IMA93_5550 : std_logic_vector(7 downto 0);
    signal IMA94_5560 : std_logic_vector(7 downto 0);
    signal IMA95_5570 : std_logic_vector(7 downto 0);
    signal IMA96_5580 : std_logic_vector(7 downto 0);
    signal IMA97_5590 : std_logic_vector(7 downto 0);
    signal IMA98_5600 : std_logic_vector(7 downto 0);
    signal IMA99_5610 : std_logic_vector(7 downto 0);
    signal IMA9_4710 : std_logic_vector(7 downto 0);
    signal IMB0_5898 : std_logic_vector(7 downto 0);
    signal IMB10_5978 : std_logic_vector(7 downto 0);
    signal IMB11_5986 : std_logic_vector(7 downto 0);
    signal IMB12_5994 : std_logic_vector(7 downto 0);
    signal IMB13_6002 : std_logic_vector(7 downto 0);
    signal IMB14_6010 : std_logic_vector(7 downto 0);
    signal IMB15_6018 : std_logic_vector(7 downto 0);
    signal IMB16_6026 : std_logic_vector(7 downto 0);
    signal IMB17_6034 : std_logic_vector(7 downto 0);
    signal IMB18_6042 : std_logic_vector(7 downto 0);
    signal IMB19_6050 : std_logic_vector(7 downto 0);
    signal IMB1_5906 : std_logic_vector(7 downto 0);
    signal IMB20_6058 : std_logic_vector(7 downto 0);
    signal IMB21_6066 : std_logic_vector(7 downto 0);
    signal IMB22_6074 : std_logic_vector(7 downto 0);
    signal IMB23_6082 : std_logic_vector(7 downto 0);
    signal IMB24_6090 : std_logic_vector(7 downto 0);
    signal IMB25_6098 : std_logic_vector(7 downto 0);
    signal IMB26_6106 : std_logic_vector(7 downto 0);
    signal IMB27_6114 : std_logic_vector(7 downto 0);
    signal IMB28_6122 : std_logic_vector(7 downto 0);
    signal IMB29_6130 : std_logic_vector(7 downto 0);
    signal IMB2_5914 : std_logic_vector(7 downto 0);
    signal IMB30_6138 : std_logic_vector(7 downto 0);
    signal IMB31_6146 : std_logic_vector(7 downto 0);
    signal IMB32_6154 : std_logic_vector(7 downto 0);
    signal IMB33_6162 : std_logic_vector(7 downto 0);
    signal IMB34_6170 : std_logic_vector(7 downto 0);
    signal IMB35_6178 : std_logic_vector(7 downto 0);
    signal IMB36_6186 : std_logic_vector(7 downto 0);
    signal IMB37_6194 : std_logic_vector(7 downto 0);
    signal IMB38_6202 : std_logic_vector(7 downto 0);
    signal IMB39_6210 : std_logic_vector(7 downto 0);
    signal IMB3_5922 : std_logic_vector(7 downto 0);
    signal IMB40_6218 : std_logic_vector(7 downto 0);
    signal IMB41_6226 : std_logic_vector(7 downto 0);
    signal IMB42_6234 : std_logic_vector(7 downto 0);
    signal IMB43_6242 : std_logic_vector(7 downto 0);
    signal IMB44_6250 : std_logic_vector(7 downto 0);
    signal IMB45_6258 : std_logic_vector(7 downto 0);
    signal IMB46_6266 : std_logic_vector(7 downto 0);
    signal IMB47_6274 : std_logic_vector(7 downto 0);
    signal IMB48_6282 : std_logic_vector(7 downto 0);
    signal IMB49_6290 : std_logic_vector(7 downto 0);
    signal IMB4_5930 : std_logic_vector(7 downto 0);
    signal IMB50_6298 : std_logic_vector(7 downto 0);
    signal IMB51_6306 : std_logic_vector(7 downto 0);
    signal IMB52_6314 : std_logic_vector(7 downto 0);
    signal IMB53_6322 : std_logic_vector(7 downto 0);
    signal IMB54_6330 : std_logic_vector(7 downto 0);
    signal IMB55_6338 : std_logic_vector(7 downto 0);
    signal IMB56_6346 : std_logic_vector(7 downto 0);
    signal IMB57_6354 : std_logic_vector(7 downto 0);
    signal IMB58_6362 : std_logic_vector(7 downto 0);
    signal IMB59_6370 : std_logic_vector(7 downto 0);
    signal IMB5_5938 : std_logic_vector(7 downto 0);
    signal IMB60_6378 : std_logic_vector(7 downto 0);
    signal IMB61_6386 : std_logic_vector(7 downto 0);
    signal IMB62_6394 : std_logic_vector(7 downto 0);
    signal IMB63_6402 : std_logic_vector(7 downto 0);
    signal IMB6_5946 : std_logic_vector(7 downto 0);
    signal IMB7_5954 : std_logic_vector(7 downto 0);
    signal IMB8_5962 : std_logic_vector(7 downto 0);
    signal IMB9_5970 : std_logic_vector(7 downto 0);
    signal IMC0_6410 : std_logic_vector(7 downto 0);
    signal IMC10_6490 : std_logic_vector(7 downto 0);
    signal IMC11_6498 : std_logic_vector(7 downto 0);
    signal IMC12_6506 : std_logic_vector(7 downto 0);
    signal IMC13_6514 : std_logic_vector(7 downto 0);
    signal IMC14_6522 : std_logic_vector(7 downto 0);
    signal IMC15_6530 : std_logic_vector(7 downto 0);
    signal IMC16_6538 : std_logic_vector(7 downto 0);
    signal IMC17_6546 : std_logic_vector(7 downto 0);
    signal IMC18_6554 : std_logic_vector(7 downto 0);
    signal IMC19_6562 : std_logic_vector(7 downto 0);
    signal IMC1_6418 : std_logic_vector(7 downto 0);
    signal IMC20_6570 : std_logic_vector(7 downto 0);
    signal IMC21_6578 : std_logic_vector(7 downto 0);
    signal IMC22_6586 : std_logic_vector(7 downto 0);
    signal IMC23_6594 : std_logic_vector(7 downto 0);
    signal IMC24_6602 : std_logic_vector(7 downto 0);
    signal IMC25_6610 : std_logic_vector(7 downto 0);
    signal IMC26_6618 : std_logic_vector(7 downto 0);
    signal IMC27_6626 : std_logic_vector(7 downto 0);
    signal IMC28_6634 : std_logic_vector(7 downto 0);
    signal IMC29_6642 : std_logic_vector(7 downto 0);
    signal IMC2_6426 : std_logic_vector(7 downto 0);
    signal IMC30_6650 : std_logic_vector(7 downto 0);
    signal IMC31_6658 : std_logic_vector(7 downto 0);
    signal IMC3_6434 : std_logic_vector(7 downto 0);
    signal IMC4_6442 : std_logic_vector(7 downto 0);
    signal IMC5_6450 : std_logic_vector(7 downto 0);
    signal IMC6_6458 : std_logic_vector(7 downto 0);
    signal IMC7_6466 : std_logic_vector(7 downto 0);
    signal IMC8_6474 : std_logic_vector(7 downto 0);
    signal IMC9_6482 : std_logic_vector(7 downto 0);
    signal IMD0_6666 : std_logic_vector(7 downto 0);
    signal IMD10_6746 : std_logic_vector(7 downto 0);
    signal IMD11_6754 : std_logic_vector(7 downto 0);
    signal IMD12_6762 : std_logic_vector(7 downto 0);
    signal IMD13_6770 : std_logic_vector(7 downto 0);
    signal IMD14_6778 : std_logic_vector(7 downto 0);
    signal IMD15_6786 : std_logic_vector(7 downto 0);
    signal IMD1_6674 : std_logic_vector(7 downto 0);
    signal IMD2_6682 : std_logic_vector(7 downto 0);
    signal IMD3_6690 : std_logic_vector(7 downto 0);
    signal IMD4_6698 : std_logic_vector(7 downto 0);
    signal IMD5_6706 : std_logic_vector(7 downto 0);
    signal IMD6_6714 : std_logic_vector(7 downto 0);
    signal IMD7_6722 : std_logic_vector(7 downto 0);
    signal IMD8_6730 : std_logic_vector(7 downto 0);
    signal IMD9_6738 : std_logic_vector(7 downto 0);
    signal IME0_6794 : std_logic_vector(7 downto 0);
    signal IME1_6802 : std_logic_vector(7 downto 0);
    signal IME2_6810 : std_logic_vector(7 downto 0);
    signal IME3_6818 : std_logic_vector(7 downto 0);
    signal IME4_6826 : std_logic_vector(7 downto 0);
    signal IME5_6834 : std_logic_vector(7 downto 0);
    signal IME6_6842 : std_logic_vector(7 downto 0);
    signal IME7_6850 : std_logic_vector(7 downto 0);
    signal IMF0_6858 : std_logic_vector(7 downto 0);
    signal IMF1_6866 : std_logic_vector(7 downto 0);
    signal IMF2_6874 : std_logic_vector(7 downto 0);
    signal IMF3_6882 : std_logic_vector(7 downto 0);
    signal IMG0_6890 : std_logic_vector(7 downto 0);
    signal IMG1_6898 : std_logic_vector(7 downto 0);
    signal konst_4613_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4623_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4633_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4643_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4653_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4663_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4673_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4683_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4693_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4703_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4713_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4723_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4733_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4743_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4753_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4763_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4773_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4783_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4793_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4803_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4813_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4823_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4833_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4843_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4853_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4863_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4873_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4883_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4893_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4903_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4913_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4923_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4933_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4943_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4953_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4963_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4973_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4983_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4993_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5003_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5013_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5023_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5033_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5043_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5053_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5063_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5073_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5083_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5093_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5103_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5113_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5123_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5133_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5143_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5153_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5163_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5173_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5183_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5193_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5203_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5213_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5223_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5233_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5243_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5253_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5263_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5273_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5283_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5293_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5303_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5313_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5323_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5333_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5343_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5353_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5363_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5373_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5383_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5393_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5403_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5413_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5423_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5433_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5443_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5453_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5463_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5473_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5483_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5493_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5503_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5513_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5523_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5533_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5543_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5553_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5563_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5573_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5583_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5593_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5603_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5613_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5623_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5633_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5643_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5653_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5663_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5673_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5683_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5693_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5703_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5713_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5723_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5733_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5743_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5753_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5763_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5773_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5783_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5793_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5803_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5813_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5823_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5833_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5843_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5853_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5863_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5873_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5883_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5893_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5901_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5909_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5917_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5925_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5933_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5941_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5949_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5957_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5965_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5973_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5981_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5989_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5997_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6005_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6013_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6021_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6029_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6037_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6045_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6053_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6061_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6069_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6077_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6085_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6093_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6101_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6109_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6117_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6125_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6133_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6141_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6149_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6157_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6165_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6173_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6181_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6189_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6197_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6205_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6213_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6221_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6229_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6237_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6245_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6253_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6261_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6269_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6277_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6285_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6293_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6301_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6309_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6317_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6325_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6333_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6341_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6349_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6357_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6365_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6373_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6381_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6389_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6397_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6405_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6413_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6421_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6429_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6437_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6445_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6453_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6461_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6469_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6477_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6485_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6493_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6501_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6509_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6517_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6525_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6533_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6541_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6549_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6557_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6565_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6573_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6581_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6589_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6597_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6605_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6613_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6621_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6629_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6637_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6645_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6653_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6661_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6669_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6677_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6685_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6693_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6701_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6709_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6717_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6725_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6733_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6741_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6749_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6757_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6765_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6773_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6781_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6789_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6797_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6805_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6813_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6821_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6829_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6837_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6845_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6853_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6861_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6869_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6877_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6885_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6893_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6901_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4616_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4618_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4626_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4628_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4636_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4638_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4646_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4648_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4656_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4658_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4666_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4668_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4676_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4678_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4686_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4688_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4696_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4698_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4706_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4708_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4716_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4718_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4726_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4728_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4736_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4738_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4746_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4748_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4756_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4758_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4766_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4768_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4776_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4778_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4786_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4788_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4796_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4798_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4806_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4808_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4816_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4818_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4826_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4828_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4836_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4838_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4846_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4848_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4856_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4858_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4866_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4868_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4876_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4878_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4886_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4888_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4896_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4898_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4906_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4908_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4916_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4918_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4926_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4928_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4936_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4938_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4946_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4948_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4956_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4958_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4966_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4968_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4976_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4978_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4986_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4988_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4996_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4998_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5006_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5008_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5016_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5018_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5026_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5028_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5036_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5038_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5046_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5048_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5056_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5058_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5066_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5068_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5076_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5078_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5086_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5088_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5096_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5098_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5106_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5108_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5116_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5118_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5126_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5128_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5136_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5138_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5146_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5148_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5156_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5158_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5166_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5168_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5176_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5178_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5186_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5188_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5196_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5198_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5206_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5208_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5216_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5218_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5226_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5228_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5236_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5238_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5246_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5248_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5256_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5258_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5266_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5268_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5276_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5278_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5286_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5288_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5296_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5298_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5306_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5308_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5316_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5318_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5326_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5328_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5336_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5338_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5346_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5348_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5356_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5358_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5366_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5368_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5376_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5378_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5386_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5388_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5396_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5398_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5406_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5408_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5416_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5418_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5426_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5428_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5436_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5438_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5446_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5448_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5456_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5458_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5466_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5468_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5476_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5478_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5486_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5488_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5496_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5498_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5506_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5508_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5516_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5518_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5526_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5528_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5536_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5538_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5546_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5548_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5556_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5558_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5566_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5568_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5576_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5578_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5586_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5588_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5596_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5598_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5606_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5608_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5616_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5618_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5626_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5628_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5636_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5638_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5646_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5648_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5656_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5658_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5666_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5668_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5676_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5678_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5686_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5688_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5696_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5698_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5706_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5708_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5716_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5718_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5726_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5728_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5736_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5738_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5746_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5748_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5756_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5758_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5766_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5768_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5776_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5778_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5786_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5788_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5796_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5798_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5806_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5808_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5816_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5818_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5826_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5828_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5836_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5838_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5846_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5848_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5856_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5858_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5866_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5868_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5876_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5878_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5886_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5888_wire_constant : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    konst_4613_wire_constant <= "00000000";
    konst_4623_wire_constant <= "00000000";
    konst_4633_wire_constant <= "00000000";
    konst_4643_wire_constant <= "00000000";
    konst_4653_wire_constant <= "00000000";
    konst_4663_wire_constant <= "00000000";
    konst_4673_wire_constant <= "00000000";
    konst_4683_wire_constant <= "00000000";
    konst_4693_wire_constant <= "00000000";
    konst_4703_wire_constant <= "00000000";
    konst_4713_wire_constant <= "00000000";
    konst_4723_wire_constant <= "00000000";
    konst_4733_wire_constant <= "00000000";
    konst_4743_wire_constant <= "00000000";
    konst_4753_wire_constant <= "00000000";
    konst_4763_wire_constant <= "00000000";
    konst_4773_wire_constant <= "00000000";
    konst_4783_wire_constant <= "00000000";
    konst_4793_wire_constant <= "00000000";
    konst_4803_wire_constant <= "00000000";
    konst_4813_wire_constant <= "00000000";
    konst_4823_wire_constant <= "00000000";
    konst_4833_wire_constant <= "00000000";
    konst_4843_wire_constant <= "00000000";
    konst_4853_wire_constant <= "00000000";
    konst_4863_wire_constant <= "00000000";
    konst_4873_wire_constant <= "00000000";
    konst_4883_wire_constant <= "00000000";
    konst_4893_wire_constant <= "00000000";
    konst_4903_wire_constant <= "00000000";
    konst_4913_wire_constant <= "00000000";
    konst_4923_wire_constant <= "00000000";
    konst_4933_wire_constant <= "00000000";
    konst_4943_wire_constant <= "00000000";
    konst_4953_wire_constant <= "00000000";
    konst_4963_wire_constant <= "00000000";
    konst_4973_wire_constant <= "00000000";
    konst_4983_wire_constant <= "00000000";
    konst_4993_wire_constant <= "00000000";
    konst_5003_wire_constant <= "00000000";
    konst_5013_wire_constant <= "00000000";
    konst_5023_wire_constant <= "00000000";
    konst_5033_wire_constant <= "00000000";
    konst_5043_wire_constant <= "00000000";
    konst_5053_wire_constant <= "00000000";
    konst_5063_wire_constant <= "00000000";
    konst_5073_wire_constant <= "00000000";
    konst_5083_wire_constant <= "00000000";
    konst_5093_wire_constant <= "00000000";
    konst_5103_wire_constant <= "00000000";
    konst_5113_wire_constant <= "00000000";
    konst_5123_wire_constant <= "00000000";
    konst_5133_wire_constant <= "00000000";
    konst_5143_wire_constant <= "00000000";
    konst_5153_wire_constant <= "00000000";
    konst_5163_wire_constant <= "00000000";
    konst_5173_wire_constant <= "00000000";
    konst_5183_wire_constant <= "00000000";
    konst_5193_wire_constant <= "00000000";
    konst_5203_wire_constant <= "00000000";
    konst_5213_wire_constant <= "00000000";
    konst_5223_wire_constant <= "00000000";
    konst_5233_wire_constant <= "00000000";
    konst_5243_wire_constant <= "00000000";
    konst_5253_wire_constant <= "00000000";
    konst_5263_wire_constant <= "00000000";
    konst_5273_wire_constant <= "00000000";
    konst_5283_wire_constant <= "00000000";
    konst_5293_wire_constant <= "00000000";
    konst_5303_wire_constant <= "00000000";
    konst_5313_wire_constant <= "00000000";
    konst_5323_wire_constant <= "00000000";
    konst_5333_wire_constant <= "00000000";
    konst_5343_wire_constant <= "00000000";
    konst_5353_wire_constant <= "00000000";
    konst_5363_wire_constant <= "00000000";
    konst_5373_wire_constant <= "00000000";
    konst_5383_wire_constant <= "00000000";
    konst_5393_wire_constant <= "00000000";
    konst_5403_wire_constant <= "00000000";
    konst_5413_wire_constant <= "00000000";
    konst_5423_wire_constant <= "00000000";
    konst_5433_wire_constant <= "00000000";
    konst_5443_wire_constant <= "00000000";
    konst_5453_wire_constant <= "00000000";
    konst_5463_wire_constant <= "00000000";
    konst_5473_wire_constant <= "00000000";
    konst_5483_wire_constant <= "00000000";
    konst_5493_wire_constant <= "00000000";
    konst_5503_wire_constant <= "00000000";
    konst_5513_wire_constant <= "00000000";
    konst_5523_wire_constant <= "00000000";
    konst_5533_wire_constant <= "00000000";
    konst_5543_wire_constant <= "00000000";
    konst_5553_wire_constant <= "00000000";
    konst_5563_wire_constant <= "00000000";
    konst_5573_wire_constant <= "00000000";
    konst_5583_wire_constant <= "00000000";
    konst_5593_wire_constant <= "00000000";
    konst_5603_wire_constant <= "00000000";
    konst_5613_wire_constant <= "00000000";
    konst_5623_wire_constant <= "00000000";
    konst_5633_wire_constant <= "00000000";
    konst_5643_wire_constant <= "00000000";
    konst_5653_wire_constant <= "00000000";
    konst_5663_wire_constant <= "00000000";
    konst_5673_wire_constant <= "00000000";
    konst_5683_wire_constant <= "00000000";
    konst_5693_wire_constant <= "00000000";
    konst_5703_wire_constant <= "00000000";
    konst_5713_wire_constant <= "00000000";
    konst_5723_wire_constant <= "00000000";
    konst_5733_wire_constant <= "00000000";
    konst_5743_wire_constant <= "00000000";
    konst_5753_wire_constant <= "00000000";
    konst_5763_wire_constant <= "00000000";
    konst_5773_wire_constant <= "00000000";
    konst_5783_wire_constant <= "00000000";
    konst_5793_wire_constant <= "00000000";
    konst_5803_wire_constant <= "00000000";
    konst_5813_wire_constant <= "00000000";
    konst_5823_wire_constant <= "00000000";
    konst_5833_wire_constant <= "00000000";
    konst_5843_wire_constant <= "00000000";
    konst_5853_wire_constant <= "00000000";
    konst_5863_wire_constant <= "00000000";
    konst_5873_wire_constant <= "00000000";
    konst_5883_wire_constant <= "00000000";
    konst_5893_wire_constant <= "00000001";
    konst_5901_wire_constant <= "00000001";
    konst_5909_wire_constant <= "00000001";
    konst_5917_wire_constant <= "00000001";
    konst_5925_wire_constant <= "00000001";
    konst_5933_wire_constant <= "00000001";
    konst_5941_wire_constant <= "00000001";
    konst_5949_wire_constant <= "00000001";
    konst_5957_wire_constant <= "00000001";
    konst_5965_wire_constant <= "00000001";
    konst_5973_wire_constant <= "00000001";
    konst_5981_wire_constant <= "00000001";
    konst_5989_wire_constant <= "00000001";
    konst_5997_wire_constant <= "00000001";
    konst_6005_wire_constant <= "00000001";
    konst_6013_wire_constant <= "00000001";
    konst_6021_wire_constant <= "00000001";
    konst_6029_wire_constant <= "00000001";
    konst_6037_wire_constant <= "00000001";
    konst_6045_wire_constant <= "00000001";
    konst_6053_wire_constant <= "00000001";
    konst_6061_wire_constant <= "00000001";
    konst_6069_wire_constant <= "00000001";
    konst_6077_wire_constant <= "00000001";
    konst_6085_wire_constant <= "00000001";
    konst_6093_wire_constant <= "00000001";
    konst_6101_wire_constant <= "00000001";
    konst_6109_wire_constant <= "00000001";
    konst_6117_wire_constant <= "00000001";
    konst_6125_wire_constant <= "00000001";
    konst_6133_wire_constant <= "00000001";
    konst_6141_wire_constant <= "00000001";
    konst_6149_wire_constant <= "00000001";
    konst_6157_wire_constant <= "00000001";
    konst_6165_wire_constant <= "00000001";
    konst_6173_wire_constant <= "00000001";
    konst_6181_wire_constant <= "00000001";
    konst_6189_wire_constant <= "00000001";
    konst_6197_wire_constant <= "00000001";
    konst_6205_wire_constant <= "00000001";
    konst_6213_wire_constant <= "00000001";
    konst_6221_wire_constant <= "00000001";
    konst_6229_wire_constant <= "00000001";
    konst_6237_wire_constant <= "00000001";
    konst_6245_wire_constant <= "00000001";
    konst_6253_wire_constant <= "00000001";
    konst_6261_wire_constant <= "00000001";
    konst_6269_wire_constant <= "00000001";
    konst_6277_wire_constant <= "00000001";
    konst_6285_wire_constant <= "00000001";
    konst_6293_wire_constant <= "00000001";
    konst_6301_wire_constant <= "00000001";
    konst_6309_wire_constant <= "00000001";
    konst_6317_wire_constant <= "00000001";
    konst_6325_wire_constant <= "00000001";
    konst_6333_wire_constant <= "00000001";
    konst_6341_wire_constant <= "00000001";
    konst_6349_wire_constant <= "00000001";
    konst_6357_wire_constant <= "00000001";
    konst_6365_wire_constant <= "00000001";
    konst_6373_wire_constant <= "00000001";
    konst_6381_wire_constant <= "00000001";
    konst_6389_wire_constant <= "00000001";
    konst_6397_wire_constant <= "00000001";
    konst_6405_wire_constant <= "00000010";
    konst_6413_wire_constant <= "00000010";
    konst_6421_wire_constant <= "00000010";
    konst_6429_wire_constant <= "00000010";
    konst_6437_wire_constant <= "00000010";
    konst_6445_wire_constant <= "00000010";
    konst_6453_wire_constant <= "00000010";
    konst_6461_wire_constant <= "00000010";
    konst_6469_wire_constant <= "00000010";
    konst_6477_wire_constant <= "00000010";
    konst_6485_wire_constant <= "00000010";
    konst_6493_wire_constant <= "00000010";
    konst_6501_wire_constant <= "00000010";
    konst_6509_wire_constant <= "00000010";
    konst_6517_wire_constant <= "00000010";
    konst_6525_wire_constant <= "00000010";
    konst_6533_wire_constant <= "00000010";
    konst_6541_wire_constant <= "00000010";
    konst_6549_wire_constant <= "00000010";
    konst_6557_wire_constant <= "00000010";
    konst_6565_wire_constant <= "00000010";
    konst_6573_wire_constant <= "00000010";
    konst_6581_wire_constant <= "00000010";
    konst_6589_wire_constant <= "00000010";
    konst_6597_wire_constant <= "00000010";
    konst_6605_wire_constant <= "00000010";
    konst_6613_wire_constant <= "00000010";
    konst_6621_wire_constant <= "00000010";
    konst_6629_wire_constant <= "00000010";
    konst_6637_wire_constant <= "00000010";
    konst_6645_wire_constant <= "00000010";
    konst_6653_wire_constant <= "00000010";
    konst_6661_wire_constant <= "00000011";
    konst_6669_wire_constant <= "00000011";
    konst_6677_wire_constant <= "00000011";
    konst_6685_wire_constant <= "00000011";
    konst_6693_wire_constant <= "00000011";
    konst_6701_wire_constant <= "00000011";
    konst_6709_wire_constant <= "00000011";
    konst_6717_wire_constant <= "00000011";
    konst_6725_wire_constant <= "00000011";
    konst_6733_wire_constant <= "00000011";
    konst_6741_wire_constant <= "00000011";
    konst_6749_wire_constant <= "00000011";
    konst_6757_wire_constant <= "00000011";
    konst_6765_wire_constant <= "00000011";
    konst_6773_wire_constant <= "00000011";
    konst_6781_wire_constant <= "00000011";
    konst_6789_wire_constant <= "00000100";
    konst_6797_wire_constant <= "00000100";
    konst_6805_wire_constant <= "00000100";
    konst_6813_wire_constant <= "00000100";
    konst_6821_wire_constant <= "00000100";
    konst_6829_wire_constant <= "00000100";
    konst_6837_wire_constant <= "00000100";
    konst_6845_wire_constant <= "00000100";
    konst_6853_wire_constant <= "00000101";
    konst_6861_wire_constant <= "00000101";
    konst_6869_wire_constant <= "00000101";
    konst_6877_wire_constant <= "00000101";
    konst_6885_wire_constant <= "00000110";
    konst_6893_wire_constant <= "00000110";
    konst_6901_wire_constant <= "00000111";
    type_cast_4616_wire_constant <= "00001001";
    type_cast_4618_wire_constant <= "01010010";
    type_cast_4626_wire_constant <= "11010101";
    type_cast_4628_wire_constant <= "01101010";
    type_cast_4636_wire_constant <= "00110110";
    type_cast_4638_wire_constant <= "00110000";
    type_cast_4646_wire_constant <= "00111000";
    type_cast_4648_wire_constant <= "10100101";
    type_cast_4656_wire_constant <= "01000000";
    type_cast_4658_wire_constant <= "10111111";
    type_cast_4666_wire_constant <= "10011110";
    type_cast_4668_wire_constant <= "10100011";
    type_cast_4676_wire_constant <= "11110011";
    type_cast_4678_wire_constant <= "10000001";
    type_cast_4686_wire_constant <= "11111011";
    type_cast_4688_wire_constant <= "11010111";
    type_cast_4696_wire_constant <= "11100011";
    type_cast_4698_wire_constant <= "01111100";
    type_cast_4706_wire_constant <= "10000010";
    type_cast_4708_wire_constant <= "00111001";
    type_cast_4716_wire_constant <= "00101111";
    type_cast_4718_wire_constant <= "10011011";
    type_cast_4726_wire_constant <= "10000111";
    type_cast_4728_wire_constant <= "11111111";
    type_cast_4736_wire_constant <= "10001110";
    type_cast_4738_wire_constant <= "00110100";
    type_cast_4746_wire_constant <= "01000100";
    type_cast_4748_wire_constant <= "01000011";
    type_cast_4756_wire_constant <= "11011110";
    type_cast_4758_wire_constant <= "11000100";
    type_cast_4766_wire_constant <= "11001011";
    type_cast_4768_wire_constant <= "11101001";
    type_cast_4776_wire_constant <= "01111011";
    type_cast_4778_wire_constant <= "01010100";
    type_cast_4786_wire_constant <= "00110010";
    type_cast_4788_wire_constant <= "10010100";
    type_cast_4796_wire_constant <= "11000010";
    type_cast_4798_wire_constant <= "10100110";
    type_cast_4806_wire_constant <= "00111101";
    type_cast_4808_wire_constant <= "00100011";
    type_cast_4816_wire_constant <= "01001100";
    type_cast_4818_wire_constant <= "11101110";
    type_cast_4826_wire_constant <= "00001011";
    type_cast_4828_wire_constant <= "10010101";
    type_cast_4836_wire_constant <= "11111010";
    type_cast_4838_wire_constant <= "01000010";
    type_cast_4846_wire_constant <= "01001110";
    type_cast_4848_wire_constant <= "11000011";
    type_cast_4856_wire_constant <= "00101110";
    type_cast_4858_wire_constant <= "00001000";
    type_cast_4866_wire_constant <= "01100110";
    type_cast_4868_wire_constant <= "10100001";
    type_cast_4876_wire_constant <= "11011001";
    type_cast_4878_wire_constant <= "00101000";
    type_cast_4886_wire_constant <= "10110010";
    type_cast_4888_wire_constant <= "00100100";
    type_cast_4896_wire_constant <= "01011011";
    type_cast_4898_wire_constant <= "01110110";
    type_cast_4906_wire_constant <= "01001001";
    type_cast_4908_wire_constant <= "10100010";
    type_cast_4916_wire_constant <= "10001011";
    type_cast_4918_wire_constant <= "01101101";
    type_cast_4926_wire_constant <= "00100101";
    type_cast_4928_wire_constant <= "11010001";
    type_cast_4936_wire_constant <= "11111000";
    type_cast_4938_wire_constant <= "01110010";
    type_cast_4946_wire_constant <= "01100100";
    type_cast_4948_wire_constant <= "11110110";
    type_cast_4956_wire_constant <= "01101000";
    type_cast_4958_wire_constant <= "10000110";
    type_cast_4966_wire_constant <= "00010110";
    type_cast_4968_wire_constant <= "10011000";
    type_cast_4976_wire_constant <= "10100100";
    type_cast_4978_wire_constant <= "11010100";
    type_cast_4986_wire_constant <= "11001100";
    type_cast_4988_wire_constant <= "01011100";
    type_cast_4996_wire_constant <= "01100101";
    type_cast_4998_wire_constant <= "01011101";
    type_cast_5006_wire_constant <= "10010010";
    type_cast_5008_wire_constant <= "10110110";
    type_cast_5016_wire_constant <= "01110000";
    type_cast_5018_wire_constant <= "01101100";
    type_cast_5026_wire_constant <= "01010000";
    type_cast_5028_wire_constant <= "01001000";
    type_cast_5036_wire_constant <= "11101101";
    type_cast_5038_wire_constant <= "11111101";
    type_cast_5046_wire_constant <= "11011010";
    type_cast_5048_wire_constant <= "10111001";
    type_cast_5056_wire_constant <= "00010101";
    type_cast_5058_wire_constant <= "01011110";
    type_cast_5066_wire_constant <= "01010111";
    type_cast_5068_wire_constant <= "01000110";
    type_cast_5076_wire_constant <= "10001101";
    type_cast_5078_wire_constant <= "10100111";
    type_cast_5086_wire_constant <= "10000100";
    type_cast_5088_wire_constant <= "10011101";
    type_cast_5096_wire_constant <= "11011000";
    type_cast_5098_wire_constant <= "10010000";
    type_cast_5106_wire_constant <= "00000000";
    type_cast_5108_wire_constant <= "10101011";
    type_cast_5116_wire_constant <= "10111100";
    type_cast_5118_wire_constant <= "10001100";
    type_cast_5126_wire_constant <= "00001010";
    type_cast_5128_wire_constant <= "11010011";
    type_cast_5136_wire_constant <= "11100100";
    type_cast_5138_wire_constant <= "11110111";
    type_cast_5146_wire_constant <= "00000101";
    type_cast_5148_wire_constant <= "01011000";
    type_cast_5156_wire_constant <= "10110011";
    type_cast_5158_wire_constant <= "10111000";
    type_cast_5166_wire_constant <= "00000110";
    type_cast_5168_wire_constant <= "01000101";
    type_cast_5176_wire_constant <= "00101100";
    type_cast_5178_wire_constant <= "11010000";
    type_cast_5186_wire_constant <= "10001111";
    type_cast_5188_wire_constant <= "00011110";
    type_cast_5196_wire_constant <= "00111111";
    type_cast_5198_wire_constant <= "11001010";
    type_cast_5206_wire_constant <= "00000010";
    type_cast_5208_wire_constant <= "00001111";
    type_cast_5216_wire_constant <= "10101111";
    type_cast_5218_wire_constant <= "11000001";
    type_cast_5226_wire_constant <= "00000011";
    type_cast_5228_wire_constant <= "10111101";
    type_cast_5236_wire_constant <= "00010011";
    type_cast_5238_wire_constant <= "00000001";
    type_cast_5246_wire_constant <= "01101011";
    type_cast_5248_wire_constant <= "10001010";
    type_cast_5256_wire_constant <= "10010001";
    type_cast_5258_wire_constant <= "00111010";
    type_cast_5266_wire_constant <= "01000001";
    type_cast_5268_wire_constant <= "00010001";
    type_cast_5276_wire_constant <= "01100111";
    type_cast_5278_wire_constant <= "01001111";
    type_cast_5286_wire_constant <= "11101010";
    type_cast_5288_wire_constant <= "11011100";
    type_cast_5296_wire_constant <= "11110010";
    type_cast_5298_wire_constant <= "10010111";
    type_cast_5306_wire_constant <= "11001110";
    type_cast_5308_wire_constant <= "11001111";
    type_cast_5316_wire_constant <= "10110100";
    type_cast_5318_wire_constant <= "11110000";
    type_cast_5326_wire_constant <= "01110011";
    type_cast_5328_wire_constant <= "11100110";
    type_cast_5336_wire_constant <= "10101100";
    type_cast_5338_wire_constant <= "10010110";
    type_cast_5346_wire_constant <= "00100010";
    type_cast_5348_wire_constant <= "01110100";
    type_cast_5356_wire_constant <= "10101101";
    type_cast_5358_wire_constant <= "11100111";
    type_cast_5366_wire_constant <= "10000101";
    type_cast_5368_wire_constant <= "00110101";
    type_cast_5376_wire_constant <= "11111001";
    type_cast_5378_wire_constant <= "11100010";
    type_cast_5386_wire_constant <= "11101000";
    type_cast_5388_wire_constant <= "00110111";
    type_cast_5396_wire_constant <= "01110101";
    type_cast_5398_wire_constant <= "00011100";
    type_cast_5406_wire_constant <= "01101110";
    type_cast_5408_wire_constant <= "11011111";
    type_cast_5416_wire_constant <= "11110001";
    type_cast_5418_wire_constant <= "01000111";
    type_cast_5426_wire_constant <= "01110001";
    type_cast_5428_wire_constant <= "00011010";
    type_cast_5436_wire_constant <= "00101001";
    type_cast_5438_wire_constant <= "00011101";
    type_cast_5446_wire_constant <= "10001001";
    type_cast_5448_wire_constant <= "11000101";
    type_cast_5456_wire_constant <= "10110111";
    type_cast_5458_wire_constant <= "01101111";
    type_cast_5466_wire_constant <= "00001110";
    type_cast_5468_wire_constant <= "01100010";
    type_cast_5476_wire_constant <= "00011000";
    type_cast_5478_wire_constant <= "10101010";
    type_cast_5486_wire_constant <= "00011011";
    type_cast_5488_wire_constant <= "10111110";
    type_cast_5496_wire_constant <= "01010110";
    type_cast_5498_wire_constant <= "11111100";
    type_cast_5506_wire_constant <= "01001011";
    type_cast_5508_wire_constant <= "00111110";
    type_cast_5516_wire_constant <= "11010010";
    type_cast_5518_wire_constant <= "11000110";
    type_cast_5526_wire_constant <= "00100000";
    type_cast_5528_wire_constant <= "01111001";
    type_cast_5536_wire_constant <= "11011011";
    type_cast_5538_wire_constant <= "10011010";
    type_cast_5546_wire_constant <= "11111110";
    type_cast_5548_wire_constant <= "11000000";
    type_cast_5556_wire_constant <= "11001101";
    type_cast_5558_wire_constant <= "01111000";
    type_cast_5566_wire_constant <= "11110100";
    type_cast_5568_wire_constant <= "01011010";
    type_cast_5576_wire_constant <= "11011101";
    type_cast_5578_wire_constant <= "00011111";
    type_cast_5586_wire_constant <= "00110011";
    type_cast_5588_wire_constant <= "10101000";
    type_cast_5596_wire_constant <= "00000111";
    type_cast_5598_wire_constant <= "10001000";
    type_cast_5606_wire_constant <= "00110001";
    type_cast_5608_wire_constant <= "11000111";
    type_cast_5616_wire_constant <= "00010010";
    type_cast_5618_wire_constant <= "10110001";
    type_cast_5626_wire_constant <= "01011001";
    type_cast_5628_wire_constant <= "00010000";
    type_cast_5636_wire_constant <= "10000000";
    type_cast_5638_wire_constant <= "00100111";
    type_cast_5646_wire_constant <= "01011111";
    type_cast_5648_wire_constant <= "11101100";
    type_cast_5656_wire_constant <= "01010001";
    type_cast_5658_wire_constant <= "01100000";
    type_cast_5666_wire_constant <= "10101001";
    type_cast_5668_wire_constant <= "01111111";
    type_cast_5676_wire_constant <= "10110101";
    type_cast_5678_wire_constant <= "00011001";
    type_cast_5686_wire_constant <= "00001101";
    type_cast_5688_wire_constant <= "01001010";
    type_cast_5696_wire_constant <= "11100101";
    type_cast_5698_wire_constant <= "00101101";
    type_cast_5706_wire_constant <= "10011111";
    type_cast_5708_wire_constant <= "01111010";
    type_cast_5716_wire_constant <= "11001001";
    type_cast_5718_wire_constant <= "10010011";
    type_cast_5726_wire_constant <= "11101111";
    type_cast_5728_wire_constant <= "10011100";
    type_cast_5736_wire_constant <= "11100000";
    type_cast_5738_wire_constant <= "10100000";
    type_cast_5746_wire_constant <= "01001101";
    type_cast_5748_wire_constant <= "00111011";
    type_cast_5756_wire_constant <= "00101010";
    type_cast_5758_wire_constant <= "10101110";
    type_cast_5766_wire_constant <= "10110000";
    type_cast_5768_wire_constant <= "11110101";
    type_cast_5776_wire_constant <= "11101011";
    type_cast_5778_wire_constant <= "11001000";
    type_cast_5786_wire_constant <= "00111100";
    type_cast_5788_wire_constant <= "10111011";
    type_cast_5796_wire_constant <= "01010011";
    type_cast_5798_wire_constant <= "10000011";
    type_cast_5806_wire_constant <= "01100001";
    type_cast_5808_wire_constant <= "10011001";
    type_cast_5816_wire_constant <= "00101011";
    type_cast_5818_wire_constant <= "00010111";
    type_cast_5826_wire_constant <= "01111110";
    type_cast_5828_wire_constant <= "00000100";
    type_cast_5836_wire_constant <= "01110111";
    type_cast_5838_wire_constant <= "10111010";
    type_cast_5846_wire_constant <= "00100110";
    type_cast_5848_wire_constant <= "11010110";
    type_cast_5856_wire_constant <= "01101001";
    type_cast_5858_wire_constant <= "11100001";
    type_cast_5866_wire_constant <= "01100011";
    type_cast_5868_wire_constant <= "00010100";
    type_cast_5876_wire_constant <= "00100001";
    type_cast_5878_wire_constant <= "01010101";
    type_cast_5886_wire_constant <= "01111101";
    type_cast_5888_wire_constant <= "00001100";
    -- logger for split-operator MUX_4619_inst flow-through 
    process(IMA0_4620) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_4619_inst:flowthrough inputs: " & " BITSEL_u8_u1_4614_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4614_wire) & " type_cast_4616_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_4616_wire_constant) & " type_cast_4618_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_4618_wire_constant) & " outputs:" & " IMA0_4620= "  & Convert_SLV_To_Hex_String(IMA0_4620));
      --
    end process; 
    -- flow-through select operator MUX_4619_inst
    IMA0_4620 <= type_cast_4616_wire_constant when (BITSEL_u8_u1_4614_wire(0) /=  '0') else type_cast_4618_wire_constant;
    -- logger for split-operator MUX_4629_inst flow-through 
    process(IMA1_4630) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_4629_inst:flowthrough inputs: " & " BITSEL_u8_u1_4624_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4624_wire) & " type_cast_4626_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_4626_wire_constant) & " type_cast_4628_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_4628_wire_constant) & " outputs:" & " IMA1_4630= "  & Convert_SLV_To_Hex_String(IMA1_4630));
      --
    end process; 
    -- flow-through select operator MUX_4629_inst
    IMA1_4630 <= type_cast_4626_wire_constant when (BITSEL_u8_u1_4624_wire(0) /=  '0') else type_cast_4628_wire_constant;
    -- logger for split-operator MUX_4639_inst flow-through 
    process(IMA2_4640) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_4639_inst:flowthrough inputs: " & " BITSEL_u8_u1_4634_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4634_wire) & " type_cast_4636_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_4636_wire_constant) & " type_cast_4638_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_4638_wire_constant) & " outputs:" & " IMA2_4640= "  & Convert_SLV_To_Hex_String(IMA2_4640));
      --
    end process; 
    -- flow-through select operator MUX_4639_inst
    IMA2_4640 <= type_cast_4636_wire_constant when (BITSEL_u8_u1_4634_wire(0) /=  '0') else type_cast_4638_wire_constant;
    -- logger for split-operator MUX_4649_inst flow-through 
    process(IMA3_4650) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_4649_inst:flowthrough inputs: " & " BITSEL_u8_u1_4644_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4644_wire) & " type_cast_4646_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_4646_wire_constant) & " type_cast_4648_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_4648_wire_constant) & " outputs:" & " IMA3_4650= "  & Convert_SLV_To_Hex_String(IMA3_4650));
      --
    end process; 
    -- flow-through select operator MUX_4649_inst
    IMA3_4650 <= type_cast_4646_wire_constant when (BITSEL_u8_u1_4644_wire(0) /=  '0') else type_cast_4648_wire_constant;
    -- logger for split-operator MUX_4659_inst flow-through 
    process(IMA4_4660) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_4659_inst:flowthrough inputs: " & " BITSEL_u8_u1_4654_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4654_wire) & " type_cast_4656_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_4656_wire_constant) & " type_cast_4658_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_4658_wire_constant) & " outputs:" & " IMA4_4660= "  & Convert_SLV_To_Hex_String(IMA4_4660));
      --
    end process; 
    -- flow-through select operator MUX_4659_inst
    IMA4_4660 <= type_cast_4656_wire_constant when (BITSEL_u8_u1_4654_wire(0) /=  '0') else type_cast_4658_wire_constant;
    -- logger for split-operator MUX_4669_inst flow-through 
    process(IMA5_4670) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_4669_inst:flowthrough inputs: " & " BITSEL_u8_u1_4664_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4664_wire) & " type_cast_4666_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_4666_wire_constant) & " type_cast_4668_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_4668_wire_constant) & " outputs:" & " IMA5_4670= "  & Convert_SLV_To_Hex_String(IMA5_4670));
      --
    end process; 
    -- flow-through select operator MUX_4669_inst
    IMA5_4670 <= type_cast_4666_wire_constant when (BITSEL_u8_u1_4664_wire(0) /=  '0') else type_cast_4668_wire_constant;
    -- logger for split-operator MUX_4679_inst flow-through 
    process(IMA6_4680) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_4679_inst:flowthrough inputs: " & " BITSEL_u8_u1_4674_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4674_wire) & " type_cast_4676_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_4676_wire_constant) & " type_cast_4678_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_4678_wire_constant) & " outputs:" & " IMA6_4680= "  & Convert_SLV_To_Hex_String(IMA6_4680));
      --
    end process; 
    -- flow-through select operator MUX_4679_inst
    IMA6_4680 <= type_cast_4676_wire_constant when (BITSEL_u8_u1_4674_wire(0) /=  '0') else type_cast_4678_wire_constant;
    -- logger for split-operator MUX_4689_inst flow-through 
    process(IMA7_4690) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_4689_inst:flowthrough inputs: " & " BITSEL_u8_u1_4684_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4684_wire) & " type_cast_4686_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_4686_wire_constant) & " type_cast_4688_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_4688_wire_constant) & " outputs:" & " IMA7_4690= "  & Convert_SLV_To_Hex_String(IMA7_4690));
      --
    end process; 
    -- flow-through select operator MUX_4689_inst
    IMA7_4690 <= type_cast_4686_wire_constant when (BITSEL_u8_u1_4684_wire(0) /=  '0') else type_cast_4688_wire_constant;
    -- logger for split-operator MUX_4699_inst flow-through 
    process(IMA8_4700) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_4699_inst:flowthrough inputs: " & " BITSEL_u8_u1_4694_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4694_wire) & " type_cast_4696_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_4696_wire_constant) & " type_cast_4698_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_4698_wire_constant) & " outputs:" & " IMA8_4700= "  & Convert_SLV_To_Hex_String(IMA8_4700));
      --
    end process; 
    -- flow-through select operator MUX_4699_inst
    IMA8_4700 <= type_cast_4696_wire_constant when (BITSEL_u8_u1_4694_wire(0) /=  '0') else type_cast_4698_wire_constant;
    -- logger for split-operator MUX_4709_inst flow-through 
    process(IMA9_4710) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_4709_inst:flowthrough inputs: " & " BITSEL_u8_u1_4704_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4704_wire) & " type_cast_4706_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_4706_wire_constant) & " type_cast_4708_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_4708_wire_constant) & " outputs:" & " IMA9_4710= "  & Convert_SLV_To_Hex_String(IMA9_4710));
      --
    end process; 
    -- flow-through select operator MUX_4709_inst
    IMA9_4710 <= type_cast_4706_wire_constant when (BITSEL_u8_u1_4704_wire(0) /=  '0') else type_cast_4708_wire_constant;
    -- logger for split-operator MUX_4719_inst flow-through 
    process(IMA10_4720) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_4719_inst:flowthrough inputs: " & " BITSEL_u8_u1_4714_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4714_wire) & " type_cast_4716_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_4716_wire_constant) & " type_cast_4718_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_4718_wire_constant) & " outputs:" & " IMA10_4720= "  & Convert_SLV_To_Hex_String(IMA10_4720));
      --
    end process; 
    -- flow-through select operator MUX_4719_inst
    IMA10_4720 <= type_cast_4716_wire_constant when (BITSEL_u8_u1_4714_wire(0) /=  '0') else type_cast_4718_wire_constant;
    -- logger for split-operator MUX_4729_inst flow-through 
    process(IMA11_4730) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_4729_inst:flowthrough inputs: " & " BITSEL_u8_u1_4724_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4724_wire) & " type_cast_4726_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_4726_wire_constant) & " type_cast_4728_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_4728_wire_constant) & " outputs:" & " IMA11_4730= "  & Convert_SLV_To_Hex_String(IMA11_4730));
      --
    end process; 
    -- flow-through select operator MUX_4729_inst
    IMA11_4730 <= type_cast_4726_wire_constant when (BITSEL_u8_u1_4724_wire(0) /=  '0') else type_cast_4728_wire_constant;
    -- logger for split-operator MUX_4739_inst flow-through 
    process(IMA12_4740) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_4739_inst:flowthrough inputs: " & " BITSEL_u8_u1_4734_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4734_wire) & " type_cast_4736_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_4736_wire_constant) & " type_cast_4738_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_4738_wire_constant) & " outputs:" & " IMA12_4740= "  & Convert_SLV_To_Hex_String(IMA12_4740));
      --
    end process; 
    -- flow-through select operator MUX_4739_inst
    IMA12_4740 <= type_cast_4736_wire_constant when (BITSEL_u8_u1_4734_wire(0) /=  '0') else type_cast_4738_wire_constant;
    -- logger for split-operator MUX_4749_inst flow-through 
    process(IMA13_4750) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_4749_inst:flowthrough inputs: " & " BITSEL_u8_u1_4744_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4744_wire) & " type_cast_4746_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_4746_wire_constant) & " type_cast_4748_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_4748_wire_constant) & " outputs:" & " IMA13_4750= "  & Convert_SLV_To_Hex_String(IMA13_4750));
      --
    end process; 
    -- flow-through select operator MUX_4749_inst
    IMA13_4750 <= type_cast_4746_wire_constant when (BITSEL_u8_u1_4744_wire(0) /=  '0') else type_cast_4748_wire_constant;
    -- logger for split-operator MUX_4759_inst flow-through 
    process(IMA14_4760) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_4759_inst:flowthrough inputs: " & " BITSEL_u8_u1_4754_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4754_wire) & " type_cast_4756_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_4756_wire_constant) & " type_cast_4758_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_4758_wire_constant) & " outputs:" & " IMA14_4760= "  & Convert_SLV_To_Hex_String(IMA14_4760));
      --
    end process; 
    -- flow-through select operator MUX_4759_inst
    IMA14_4760 <= type_cast_4756_wire_constant when (BITSEL_u8_u1_4754_wire(0) /=  '0') else type_cast_4758_wire_constant;
    -- logger for split-operator MUX_4769_inst flow-through 
    process(IMA15_4770) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_4769_inst:flowthrough inputs: " & " BITSEL_u8_u1_4764_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4764_wire) & " type_cast_4766_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_4766_wire_constant) & " type_cast_4768_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_4768_wire_constant) & " outputs:" & " IMA15_4770= "  & Convert_SLV_To_Hex_String(IMA15_4770));
      --
    end process; 
    -- flow-through select operator MUX_4769_inst
    IMA15_4770 <= type_cast_4766_wire_constant when (BITSEL_u8_u1_4764_wire(0) /=  '0') else type_cast_4768_wire_constant;
    -- logger for split-operator MUX_4779_inst flow-through 
    process(IMA16_4780) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_4779_inst:flowthrough inputs: " & " BITSEL_u8_u1_4774_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4774_wire) & " type_cast_4776_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_4776_wire_constant) & " type_cast_4778_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_4778_wire_constant) & " outputs:" & " IMA16_4780= "  & Convert_SLV_To_Hex_String(IMA16_4780));
      --
    end process; 
    -- flow-through select operator MUX_4779_inst
    IMA16_4780 <= type_cast_4776_wire_constant when (BITSEL_u8_u1_4774_wire(0) /=  '0') else type_cast_4778_wire_constant;
    -- logger for split-operator MUX_4789_inst flow-through 
    process(IMA17_4790) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_4789_inst:flowthrough inputs: " & " BITSEL_u8_u1_4784_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4784_wire) & " type_cast_4786_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_4786_wire_constant) & " type_cast_4788_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_4788_wire_constant) & " outputs:" & " IMA17_4790= "  & Convert_SLV_To_Hex_String(IMA17_4790));
      --
    end process; 
    -- flow-through select operator MUX_4789_inst
    IMA17_4790 <= type_cast_4786_wire_constant when (BITSEL_u8_u1_4784_wire(0) /=  '0') else type_cast_4788_wire_constant;
    -- logger for split-operator MUX_4799_inst flow-through 
    process(IMA18_4800) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_4799_inst:flowthrough inputs: " & " BITSEL_u8_u1_4794_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4794_wire) & " type_cast_4796_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_4796_wire_constant) & " type_cast_4798_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_4798_wire_constant) & " outputs:" & " IMA18_4800= "  & Convert_SLV_To_Hex_String(IMA18_4800));
      --
    end process; 
    -- flow-through select operator MUX_4799_inst
    IMA18_4800 <= type_cast_4796_wire_constant when (BITSEL_u8_u1_4794_wire(0) /=  '0') else type_cast_4798_wire_constant;
    -- logger for split-operator MUX_4809_inst flow-through 
    process(IMA19_4810) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_4809_inst:flowthrough inputs: " & " BITSEL_u8_u1_4804_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4804_wire) & " type_cast_4806_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_4806_wire_constant) & " type_cast_4808_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_4808_wire_constant) & " outputs:" & " IMA19_4810= "  & Convert_SLV_To_Hex_String(IMA19_4810));
      --
    end process; 
    -- flow-through select operator MUX_4809_inst
    IMA19_4810 <= type_cast_4806_wire_constant when (BITSEL_u8_u1_4804_wire(0) /=  '0') else type_cast_4808_wire_constant;
    -- logger for split-operator MUX_4819_inst flow-through 
    process(IMA20_4820) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_4819_inst:flowthrough inputs: " & " BITSEL_u8_u1_4814_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4814_wire) & " type_cast_4816_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_4816_wire_constant) & " type_cast_4818_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_4818_wire_constant) & " outputs:" & " IMA20_4820= "  & Convert_SLV_To_Hex_String(IMA20_4820));
      --
    end process; 
    -- flow-through select operator MUX_4819_inst
    IMA20_4820 <= type_cast_4816_wire_constant when (BITSEL_u8_u1_4814_wire(0) /=  '0') else type_cast_4818_wire_constant;
    -- logger for split-operator MUX_4829_inst flow-through 
    process(IMA21_4830) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_4829_inst:flowthrough inputs: " & " BITSEL_u8_u1_4824_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4824_wire) & " type_cast_4826_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_4826_wire_constant) & " type_cast_4828_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_4828_wire_constant) & " outputs:" & " IMA21_4830= "  & Convert_SLV_To_Hex_String(IMA21_4830));
      --
    end process; 
    -- flow-through select operator MUX_4829_inst
    IMA21_4830 <= type_cast_4826_wire_constant when (BITSEL_u8_u1_4824_wire(0) /=  '0') else type_cast_4828_wire_constant;
    -- logger for split-operator MUX_4839_inst flow-through 
    process(IMA22_4840) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_4839_inst:flowthrough inputs: " & " BITSEL_u8_u1_4834_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4834_wire) & " type_cast_4836_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_4836_wire_constant) & " type_cast_4838_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_4838_wire_constant) & " outputs:" & " IMA22_4840= "  & Convert_SLV_To_Hex_String(IMA22_4840));
      --
    end process; 
    -- flow-through select operator MUX_4839_inst
    IMA22_4840 <= type_cast_4836_wire_constant when (BITSEL_u8_u1_4834_wire(0) /=  '0') else type_cast_4838_wire_constant;
    -- logger for split-operator MUX_4849_inst flow-through 
    process(IMA23_4850) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_4849_inst:flowthrough inputs: " & " BITSEL_u8_u1_4844_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4844_wire) & " type_cast_4846_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_4846_wire_constant) & " type_cast_4848_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_4848_wire_constant) & " outputs:" & " IMA23_4850= "  & Convert_SLV_To_Hex_String(IMA23_4850));
      --
    end process; 
    -- flow-through select operator MUX_4849_inst
    IMA23_4850 <= type_cast_4846_wire_constant when (BITSEL_u8_u1_4844_wire(0) /=  '0') else type_cast_4848_wire_constant;
    -- logger for split-operator MUX_4859_inst flow-through 
    process(IMA24_4860) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_4859_inst:flowthrough inputs: " & " BITSEL_u8_u1_4854_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4854_wire) & " type_cast_4856_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_4856_wire_constant) & " type_cast_4858_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_4858_wire_constant) & " outputs:" & " IMA24_4860= "  & Convert_SLV_To_Hex_String(IMA24_4860));
      --
    end process; 
    -- flow-through select operator MUX_4859_inst
    IMA24_4860 <= type_cast_4856_wire_constant when (BITSEL_u8_u1_4854_wire(0) /=  '0') else type_cast_4858_wire_constant;
    -- logger for split-operator MUX_4869_inst flow-through 
    process(IMA25_4870) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_4869_inst:flowthrough inputs: " & " BITSEL_u8_u1_4864_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4864_wire) & " type_cast_4866_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_4866_wire_constant) & " type_cast_4868_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_4868_wire_constant) & " outputs:" & " IMA25_4870= "  & Convert_SLV_To_Hex_String(IMA25_4870));
      --
    end process; 
    -- flow-through select operator MUX_4869_inst
    IMA25_4870 <= type_cast_4866_wire_constant when (BITSEL_u8_u1_4864_wire(0) /=  '0') else type_cast_4868_wire_constant;
    -- logger for split-operator MUX_4879_inst flow-through 
    process(IMA26_4880) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_4879_inst:flowthrough inputs: " & " BITSEL_u8_u1_4874_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4874_wire) & " type_cast_4876_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_4876_wire_constant) & " type_cast_4878_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_4878_wire_constant) & " outputs:" & " IMA26_4880= "  & Convert_SLV_To_Hex_String(IMA26_4880));
      --
    end process; 
    -- flow-through select operator MUX_4879_inst
    IMA26_4880 <= type_cast_4876_wire_constant when (BITSEL_u8_u1_4874_wire(0) /=  '0') else type_cast_4878_wire_constant;
    -- logger for split-operator MUX_4889_inst flow-through 
    process(IMA27_4890) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_4889_inst:flowthrough inputs: " & " BITSEL_u8_u1_4884_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4884_wire) & " type_cast_4886_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_4886_wire_constant) & " type_cast_4888_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_4888_wire_constant) & " outputs:" & " IMA27_4890= "  & Convert_SLV_To_Hex_String(IMA27_4890));
      --
    end process; 
    -- flow-through select operator MUX_4889_inst
    IMA27_4890 <= type_cast_4886_wire_constant when (BITSEL_u8_u1_4884_wire(0) /=  '0') else type_cast_4888_wire_constant;
    -- logger for split-operator MUX_4899_inst flow-through 
    process(IMA28_4900) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_4899_inst:flowthrough inputs: " & " BITSEL_u8_u1_4894_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4894_wire) & " type_cast_4896_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_4896_wire_constant) & " type_cast_4898_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_4898_wire_constant) & " outputs:" & " IMA28_4900= "  & Convert_SLV_To_Hex_String(IMA28_4900));
      --
    end process; 
    -- flow-through select operator MUX_4899_inst
    IMA28_4900 <= type_cast_4896_wire_constant when (BITSEL_u8_u1_4894_wire(0) /=  '0') else type_cast_4898_wire_constant;
    -- logger for split-operator MUX_4909_inst flow-through 
    process(IMA29_4910) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_4909_inst:flowthrough inputs: " & " BITSEL_u8_u1_4904_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4904_wire) & " type_cast_4906_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_4906_wire_constant) & " type_cast_4908_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_4908_wire_constant) & " outputs:" & " IMA29_4910= "  & Convert_SLV_To_Hex_String(IMA29_4910));
      --
    end process; 
    -- flow-through select operator MUX_4909_inst
    IMA29_4910 <= type_cast_4906_wire_constant when (BITSEL_u8_u1_4904_wire(0) /=  '0') else type_cast_4908_wire_constant;
    -- logger for split-operator MUX_4919_inst flow-through 
    process(IMA30_4920) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_4919_inst:flowthrough inputs: " & " BITSEL_u8_u1_4914_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4914_wire) & " type_cast_4916_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_4916_wire_constant) & " type_cast_4918_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_4918_wire_constant) & " outputs:" & " IMA30_4920= "  & Convert_SLV_To_Hex_String(IMA30_4920));
      --
    end process; 
    -- flow-through select operator MUX_4919_inst
    IMA30_4920 <= type_cast_4916_wire_constant when (BITSEL_u8_u1_4914_wire(0) /=  '0') else type_cast_4918_wire_constant;
    -- logger for split-operator MUX_4929_inst flow-through 
    process(IMA31_4930) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_4929_inst:flowthrough inputs: " & " BITSEL_u8_u1_4924_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4924_wire) & " type_cast_4926_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_4926_wire_constant) & " type_cast_4928_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_4928_wire_constant) & " outputs:" & " IMA31_4930= "  & Convert_SLV_To_Hex_String(IMA31_4930));
      --
    end process; 
    -- flow-through select operator MUX_4929_inst
    IMA31_4930 <= type_cast_4926_wire_constant when (BITSEL_u8_u1_4924_wire(0) /=  '0') else type_cast_4928_wire_constant;
    -- logger for split-operator MUX_4939_inst flow-through 
    process(IMA32_4940) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_4939_inst:flowthrough inputs: " & " BITSEL_u8_u1_4934_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4934_wire) & " type_cast_4936_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_4936_wire_constant) & " type_cast_4938_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_4938_wire_constant) & " outputs:" & " IMA32_4940= "  & Convert_SLV_To_Hex_String(IMA32_4940));
      --
    end process; 
    -- flow-through select operator MUX_4939_inst
    IMA32_4940 <= type_cast_4936_wire_constant when (BITSEL_u8_u1_4934_wire(0) /=  '0') else type_cast_4938_wire_constant;
    -- logger for split-operator MUX_4949_inst flow-through 
    process(IMA33_4950) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_4949_inst:flowthrough inputs: " & " BITSEL_u8_u1_4944_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4944_wire) & " type_cast_4946_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_4946_wire_constant) & " type_cast_4948_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_4948_wire_constant) & " outputs:" & " IMA33_4950= "  & Convert_SLV_To_Hex_String(IMA33_4950));
      --
    end process; 
    -- flow-through select operator MUX_4949_inst
    IMA33_4950 <= type_cast_4946_wire_constant when (BITSEL_u8_u1_4944_wire(0) /=  '0') else type_cast_4948_wire_constant;
    -- logger for split-operator MUX_4959_inst flow-through 
    process(IMA34_4960) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_4959_inst:flowthrough inputs: " & " BITSEL_u8_u1_4954_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4954_wire) & " type_cast_4956_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_4956_wire_constant) & " type_cast_4958_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_4958_wire_constant) & " outputs:" & " IMA34_4960= "  & Convert_SLV_To_Hex_String(IMA34_4960));
      --
    end process; 
    -- flow-through select operator MUX_4959_inst
    IMA34_4960 <= type_cast_4956_wire_constant when (BITSEL_u8_u1_4954_wire(0) /=  '0') else type_cast_4958_wire_constant;
    -- logger for split-operator MUX_4969_inst flow-through 
    process(IMA35_4970) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_4969_inst:flowthrough inputs: " & " BITSEL_u8_u1_4964_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4964_wire) & " type_cast_4966_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_4966_wire_constant) & " type_cast_4968_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_4968_wire_constant) & " outputs:" & " IMA35_4970= "  & Convert_SLV_To_Hex_String(IMA35_4970));
      --
    end process; 
    -- flow-through select operator MUX_4969_inst
    IMA35_4970 <= type_cast_4966_wire_constant when (BITSEL_u8_u1_4964_wire(0) /=  '0') else type_cast_4968_wire_constant;
    -- logger for split-operator MUX_4979_inst flow-through 
    process(IMA36_4980) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_4979_inst:flowthrough inputs: " & " BITSEL_u8_u1_4974_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4974_wire) & " type_cast_4976_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_4976_wire_constant) & " type_cast_4978_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_4978_wire_constant) & " outputs:" & " IMA36_4980= "  & Convert_SLV_To_Hex_String(IMA36_4980));
      --
    end process; 
    -- flow-through select operator MUX_4979_inst
    IMA36_4980 <= type_cast_4976_wire_constant when (BITSEL_u8_u1_4974_wire(0) /=  '0') else type_cast_4978_wire_constant;
    -- logger for split-operator MUX_4989_inst flow-through 
    process(IMA37_4990) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_4989_inst:flowthrough inputs: " & " BITSEL_u8_u1_4984_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4984_wire) & " type_cast_4986_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_4986_wire_constant) & " type_cast_4988_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_4988_wire_constant) & " outputs:" & " IMA37_4990= "  & Convert_SLV_To_Hex_String(IMA37_4990));
      --
    end process; 
    -- flow-through select operator MUX_4989_inst
    IMA37_4990 <= type_cast_4986_wire_constant when (BITSEL_u8_u1_4984_wire(0) /=  '0') else type_cast_4988_wire_constant;
    -- logger for split-operator MUX_4999_inst flow-through 
    process(IMA38_5000) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_4999_inst:flowthrough inputs: " & " BITSEL_u8_u1_4994_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_4994_wire) & " type_cast_4996_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_4996_wire_constant) & " type_cast_4998_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_4998_wire_constant) & " outputs:" & " IMA38_5000= "  & Convert_SLV_To_Hex_String(IMA38_5000));
      --
    end process; 
    -- flow-through select operator MUX_4999_inst
    IMA38_5000 <= type_cast_4996_wire_constant when (BITSEL_u8_u1_4994_wire(0) /=  '0') else type_cast_4998_wire_constant;
    -- logger for split-operator MUX_5009_inst flow-through 
    process(IMA39_5010) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_5009_inst:flowthrough inputs: " & " BITSEL_u8_u1_5004_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_5004_wire) & " type_cast_5006_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5006_wire_constant) & " type_cast_5008_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5008_wire_constant) & " outputs:" & " IMA39_5010= "  & Convert_SLV_To_Hex_String(IMA39_5010));
      --
    end process; 
    -- flow-through select operator MUX_5009_inst
    IMA39_5010 <= type_cast_5006_wire_constant when (BITSEL_u8_u1_5004_wire(0) /=  '0') else type_cast_5008_wire_constant;
    -- logger for split-operator MUX_5019_inst flow-through 
    process(IMA40_5020) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_5019_inst:flowthrough inputs: " & " BITSEL_u8_u1_5014_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_5014_wire) & " type_cast_5016_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5016_wire_constant) & " type_cast_5018_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5018_wire_constant) & " outputs:" & " IMA40_5020= "  & Convert_SLV_To_Hex_String(IMA40_5020));
      --
    end process; 
    -- flow-through select operator MUX_5019_inst
    IMA40_5020 <= type_cast_5016_wire_constant when (BITSEL_u8_u1_5014_wire(0) /=  '0') else type_cast_5018_wire_constant;
    -- logger for split-operator MUX_5029_inst flow-through 
    process(IMA41_5030) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_5029_inst:flowthrough inputs: " & " BITSEL_u8_u1_5024_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_5024_wire) & " type_cast_5026_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5026_wire_constant) & " type_cast_5028_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5028_wire_constant) & " outputs:" & " IMA41_5030= "  & Convert_SLV_To_Hex_String(IMA41_5030));
      --
    end process; 
    -- flow-through select operator MUX_5029_inst
    IMA41_5030 <= type_cast_5026_wire_constant when (BITSEL_u8_u1_5024_wire(0) /=  '0') else type_cast_5028_wire_constant;
    -- logger for split-operator MUX_5039_inst flow-through 
    process(IMA42_5040) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_5039_inst:flowthrough inputs: " & " BITSEL_u8_u1_5034_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_5034_wire) & " type_cast_5036_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5036_wire_constant) & " type_cast_5038_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5038_wire_constant) & " outputs:" & " IMA42_5040= "  & Convert_SLV_To_Hex_String(IMA42_5040));
      --
    end process; 
    -- flow-through select operator MUX_5039_inst
    IMA42_5040 <= type_cast_5036_wire_constant when (BITSEL_u8_u1_5034_wire(0) /=  '0') else type_cast_5038_wire_constant;
    -- logger for split-operator MUX_5049_inst flow-through 
    process(IMA43_5050) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_5049_inst:flowthrough inputs: " & " BITSEL_u8_u1_5044_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_5044_wire) & " type_cast_5046_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5046_wire_constant) & " type_cast_5048_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5048_wire_constant) & " outputs:" & " IMA43_5050= "  & Convert_SLV_To_Hex_String(IMA43_5050));
      --
    end process; 
    -- flow-through select operator MUX_5049_inst
    IMA43_5050 <= type_cast_5046_wire_constant when (BITSEL_u8_u1_5044_wire(0) /=  '0') else type_cast_5048_wire_constant;
    -- logger for split-operator MUX_5059_inst flow-through 
    process(IMA44_5060) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_5059_inst:flowthrough inputs: " & " BITSEL_u8_u1_5054_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_5054_wire) & " type_cast_5056_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5056_wire_constant) & " type_cast_5058_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5058_wire_constant) & " outputs:" & " IMA44_5060= "  & Convert_SLV_To_Hex_String(IMA44_5060));
      --
    end process; 
    -- flow-through select operator MUX_5059_inst
    IMA44_5060 <= type_cast_5056_wire_constant when (BITSEL_u8_u1_5054_wire(0) /=  '0') else type_cast_5058_wire_constant;
    -- logger for split-operator MUX_5069_inst flow-through 
    process(IMA45_5070) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_5069_inst:flowthrough inputs: " & " BITSEL_u8_u1_5064_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_5064_wire) & " type_cast_5066_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5066_wire_constant) & " type_cast_5068_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5068_wire_constant) & " outputs:" & " IMA45_5070= "  & Convert_SLV_To_Hex_String(IMA45_5070));
      --
    end process; 
    -- flow-through select operator MUX_5069_inst
    IMA45_5070 <= type_cast_5066_wire_constant when (BITSEL_u8_u1_5064_wire(0) /=  '0') else type_cast_5068_wire_constant;
    -- logger for split-operator MUX_5079_inst flow-through 
    process(IMA46_5080) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_5079_inst:flowthrough inputs: " & " BITSEL_u8_u1_5074_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_5074_wire) & " type_cast_5076_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5076_wire_constant) & " type_cast_5078_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5078_wire_constant) & " outputs:" & " IMA46_5080= "  & Convert_SLV_To_Hex_String(IMA46_5080));
      --
    end process; 
    -- flow-through select operator MUX_5079_inst
    IMA46_5080 <= type_cast_5076_wire_constant when (BITSEL_u8_u1_5074_wire(0) /=  '0') else type_cast_5078_wire_constant;
    -- logger for split-operator MUX_5089_inst flow-through 
    process(IMA47_5090) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_5089_inst:flowthrough inputs: " & " BITSEL_u8_u1_5084_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_5084_wire) & " type_cast_5086_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5086_wire_constant) & " type_cast_5088_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5088_wire_constant) & " outputs:" & " IMA47_5090= "  & Convert_SLV_To_Hex_String(IMA47_5090));
      --
    end process; 
    -- flow-through select operator MUX_5089_inst
    IMA47_5090 <= type_cast_5086_wire_constant when (BITSEL_u8_u1_5084_wire(0) /=  '0') else type_cast_5088_wire_constant;
    -- logger for split-operator MUX_5099_inst flow-through 
    process(IMA48_5100) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_5099_inst:flowthrough inputs: " & " BITSEL_u8_u1_5094_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_5094_wire) & " type_cast_5096_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5096_wire_constant) & " type_cast_5098_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5098_wire_constant) & " outputs:" & " IMA48_5100= "  & Convert_SLV_To_Hex_String(IMA48_5100));
      --
    end process; 
    -- flow-through select operator MUX_5099_inst
    IMA48_5100 <= type_cast_5096_wire_constant when (BITSEL_u8_u1_5094_wire(0) /=  '0') else type_cast_5098_wire_constant;
    -- logger for split-operator MUX_5109_inst flow-through 
    process(IMA49_5110) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_5109_inst:flowthrough inputs: " & " BITSEL_u8_u1_5104_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_5104_wire) & " type_cast_5106_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5106_wire_constant) & " type_cast_5108_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5108_wire_constant) & " outputs:" & " IMA49_5110= "  & Convert_SLV_To_Hex_String(IMA49_5110));
      --
    end process; 
    -- flow-through select operator MUX_5109_inst
    IMA49_5110 <= type_cast_5106_wire_constant when (BITSEL_u8_u1_5104_wire(0) /=  '0') else type_cast_5108_wire_constant;
    -- logger for split-operator MUX_5119_inst flow-through 
    process(IMA50_5120) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_5119_inst:flowthrough inputs: " & " BITSEL_u8_u1_5114_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_5114_wire) & " type_cast_5116_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5116_wire_constant) & " type_cast_5118_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5118_wire_constant) & " outputs:" & " IMA50_5120= "  & Convert_SLV_To_Hex_String(IMA50_5120));
      --
    end process; 
    -- flow-through select operator MUX_5119_inst
    IMA50_5120 <= type_cast_5116_wire_constant when (BITSEL_u8_u1_5114_wire(0) /=  '0') else type_cast_5118_wire_constant;
    -- logger for split-operator MUX_5129_inst flow-through 
    process(IMA51_5130) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_5129_inst:flowthrough inputs: " & " BITSEL_u8_u1_5124_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_5124_wire) & " type_cast_5126_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5126_wire_constant) & " type_cast_5128_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5128_wire_constant) & " outputs:" & " IMA51_5130= "  & Convert_SLV_To_Hex_String(IMA51_5130));
      --
    end process; 
    -- flow-through select operator MUX_5129_inst
    IMA51_5130 <= type_cast_5126_wire_constant when (BITSEL_u8_u1_5124_wire(0) /=  '0') else type_cast_5128_wire_constant;
    -- logger for split-operator MUX_5139_inst flow-through 
    process(IMA52_5140) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_5139_inst:flowthrough inputs: " & " BITSEL_u8_u1_5134_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_5134_wire) & " type_cast_5136_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5136_wire_constant) & " type_cast_5138_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5138_wire_constant) & " outputs:" & " IMA52_5140= "  & Convert_SLV_To_Hex_String(IMA52_5140));
      --
    end process; 
    -- flow-through select operator MUX_5139_inst
    IMA52_5140 <= type_cast_5136_wire_constant when (BITSEL_u8_u1_5134_wire(0) /=  '0') else type_cast_5138_wire_constant;
    -- logger for split-operator MUX_5149_inst flow-through 
    process(IMA53_5150) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_5149_inst:flowthrough inputs: " & " BITSEL_u8_u1_5144_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_5144_wire) & " type_cast_5146_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5146_wire_constant) & " type_cast_5148_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5148_wire_constant) & " outputs:" & " IMA53_5150= "  & Convert_SLV_To_Hex_String(IMA53_5150));
      --
    end process; 
    -- flow-through select operator MUX_5149_inst
    IMA53_5150 <= type_cast_5146_wire_constant when (BITSEL_u8_u1_5144_wire(0) /=  '0') else type_cast_5148_wire_constant;
    -- logger for split-operator MUX_5159_inst flow-through 
    process(IMA54_5160) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_5159_inst:flowthrough inputs: " & " BITSEL_u8_u1_5154_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_5154_wire) & " type_cast_5156_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5156_wire_constant) & " type_cast_5158_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5158_wire_constant) & " outputs:" & " IMA54_5160= "  & Convert_SLV_To_Hex_String(IMA54_5160));
      --
    end process; 
    -- flow-through select operator MUX_5159_inst
    IMA54_5160 <= type_cast_5156_wire_constant when (BITSEL_u8_u1_5154_wire(0) /=  '0') else type_cast_5158_wire_constant;
    -- logger for split-operator MUX_5169_inst flow-through 
    process(IMA55_5170) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_5169_inst:flowthrough inputs: " & " BITSEL_u8_u1_5164_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_5164_wire) & " type_cast_5166_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5166_wire_constant) & " type_cast_5168_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5168_wire_constant) & " outputs:" & " IMA55_5170= "  & Convert_SLV_To_Hex_String(IMA55_5170));
      --
    end process; 
    -- flow-through select operator MUX_5169_inst
    IMA55_5170 <= type_cast_5166_wire_constant when (BITSEL_u8_u1_5164_wire(0) /=  '0') else type_cast_5168_wire_constant;
    -- logger for split-operator MUX_5179_inst flow-through 
    process(IMA56_5180) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_5179_inst:flowthrough inputs: " & " BITSEL_u8_u1_5174_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_5174_wire) & " type_cast_5176_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5176_wire_constant) & " type_cast_5178_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5178_wire_constant) & " outputs:" & " IMA56_5180= "  & Convert_SLV_To_Hex_String(IMA56_5180));
      --
    end process; 
    -- flow-through select operator MUX_5179_inst
    IMA56_5180 <= type_cast_5176_wire_constant when (BITSEL_u8_u1_5174_wire(0) /=  '0') else type_cast_5178_wire_constant;
    -- logger for split-operator MUX_5189_inst flow-through 
    process(IMA57_5190) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_5189_inst:flowthrough inputs: " & " BITSEL_u8_u1_5184_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_5184_wire) & " type_cast_5186_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5186_wire_constant) & " type_cast_5188_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5188_wire_constant) & " outputs:" & " IMA57_5190= "  & Convert_SLV_To_Hex_String(IMA57_5190));
      --
    end process; 
    -- flow-through select operator MUX_5189_inst
    IMA57_5190 <= type_cast_5186_wire_constant when (BITSEL_u8_u1_5184_wire(0) /=  '0') else type_cast_5188_wire_constant;
    -- logger for split-operator MUX_5199_inst flow-through 
    process(IMA58_5200) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_5199_inst:flowthrough inputs: " & " BITSEL_u8_u1_5194_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_5194_wire) & " type_cast_5196_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5196_wire_constant) & " type_cast_5198_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5198_wire_constant) & " outputs:" & " IMA58_5200= "  & Convert_SLV_To_Hex_String(IMA58_5200));
      --
    end process; 
    -- flow-through select operator MUX_5199_inst
    IMA58_5200 <= type_cast_5196_wire_constant when (BITSEL_u8_u1_5194_wire(0) /=  '0') else type_cast_5198_wire_constant;
    -- logger for split-operator MUX_5209_inst flow-through 
    process(IMA59_5210) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_5209_inst:flowthrough inputs: " & " BITSEL_u8_u1_5204_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_5204_wire) & " type_cast_5206_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5206_wire_constant) & " type_cast_5208_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5208_wire_constant) & " outputs:" & " IMA59_5210= "  & Convert_SLV_To_Hex_String(IMA59_5210));
      --
    end process; 
    -- flow-through select operator MUX_5209_inst
    IMA59_5210 <= type_cast_5206_wire_constant when (BITSEL_u8_u1_5204_wire(0) /=  '0') else type_cast_5208_wire_constant;
    -- logger for split-operator MUX_5219_inst flow-through 
    process(IMA60_5220) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_5219_inst:flowthrough inputs: " & " BITSEL_u8_u1_5214_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_5214_wire) & " type_cast_5216_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5216_wire_constant) & " type_cast_5218_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5218_wire_constant) & " outputs:" & " IMA60_5220= "  & Convert_SLV_To_Hex_String(IMA60_5220));
      --
    end process; 
    -- flow-through select operator MUX_5219_inst
    IMA60_5220 <= type_cast_5216_wire_constant when (BITSEL_u8_u1_5214_wire(0) /=  '0') else type_cast_5218_wire_constant;
    -- logger for split-operator MUX_5229_inst flow-through 
    process(IMA61_5230) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_5229_inst:flowthrough inputs: " & " BITSEL_u8_u1_5224_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_5224_wire) & " type_cast_5226_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5226_wire_constant) & " type_cast_5228_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5228_wire_constant) & " outputs:" & " IMA61_5230= "  & Convert_SLV_To_Hex_String(IMA61_5230));
      --
    end process; 
    -- flow-through select operator MUX_5229_inst
    IMA61_5230 <= type_cast_5226_wire_constant when (BITSEL_u8_u1_5224_wire(0) /=  '0') else type_cast_5228_wire_constant;
    -- logger for split-operator MUX_5239_inst flow-through 
    process(IMA62_5240) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_5239_inst:flowthrough inputs: " & " BITSEL_u8_u1_5234_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_5234_wire) & " type_cast_5236_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5236_wire_constant) & " type_cast_5238_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5238_wire_constant) & " outputs:" & " IMA62_5240= "  & Convert_SLV_To_Hex_String(IMA62_5240));
      --
    end process; 
    -- flow-through select operator MUX_5239_inst
    IMA62_5240 <= type_cast_5236_wire_constant when (BITSEL_u8_u1_5234_wire(0) /=  '0') else type_cast_5238_wire_constant;
    -- logger for split-operator MUX_5249_inst flow-through 
    process(IMA63_5250) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_5249_inst:flowthrough inputs: " & " BITSEL_u8_u1_5244_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_5244_wire) & " type_cast_5246_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5246_wire_constant) & " type_cast_5248_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5248_wire_constant) & " outputs:" & " IMA63_5250= "  & Convert_SLV_To_Hex_String(IMA63_5250));
      --
    end process; 
    -- flow-through select operator MUX_5249_inst
    IMA63_5250 <= type_cast_5246_wire_constant when (BITSEL_u8_u1_5244_wire(0) /=  '0') else type_cast_5248_wire_constant;
    -- logger for split-operator MUX_5259_inst flow-through 
    process(IMA64_5260) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_5259_inst:flowthrough inputs: " & " BITSEL_u8_u1_5254_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_5254_wire) & " type_cast_5256_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5256_wire_constant) & " type_cast_5258_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5258_wire_constant) & " outputs:" & " IMA64_5260= "  & Convert_SLV_To_Hex_String(IMA64_5260));
      --
    end process; 
    -- flow-through select operator MUX_5259_inst
    IMA64_5260 <= type_cast_5256_wire_constant when (BITSEL_u8_u1_5254_wire(0) /=  '0') else type_cast_5258_wire_constant;
    -- logger for split-operator MUX_5269_inst flow-through 
    process(IMA65_5270) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_5269_inst:flowthrough inputs: " & " BITSEL_u8_u1_5264_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_5264_wire) & " type_cast_5266_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5266_wire_constant) & " type_cast_5268_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5268_wire_constant) & " outputs:" & " IMA65_5270= "  & Convert_SLV_To_Hex_String(IMA65_5270));
      --
    end process; 
    -- flow-through select operator MUX_5269_inst
    IMA65_5270 <= type_cast_5266_wire_constant when (BITSEL_u8_u1_5264_wire(0) /=  '0') else type_cast_5268_wire_constant;
    -- logger for split-operator MUX_5279_inst flow-through 
    process(IMA66_5280) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_5279_inst:flowthrough inputs: " & " BITSEL_u8_u1_5274_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_5274_wire) & " type_cast_5276_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5276_wire_constant) & " type_cast_5278_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5278_wire_constant) & " outputs:" & " IMA66_5280= "  & Convert_SLV_To_Hex_String(IMA66_5280));
      --
    end process; 
    -- flow-through select operator MUX_5279_inst
    IMA66_5280 <= type_cast_5276_wire_constant when (BITSEL_u8_u1_5274_wire(0) /=  '0') else type_cast_5278_wire_constant;
    -- logger for split-operator MUX_5289_inst flow-through 
    process(IMA67_5290) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_5289_inst:flowthrough inputs: " & " BITSEL_u8_u1_5284_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_5284_wire) & " type_cast_5286_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5286_wire_constant) & " type_cast_5288_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5288_wire_constant) & " outputs:" & " IMA67_5290= "  & Convert_SLV_To_Hex_String(IMA67_5290));
      --
    end process; 
    -- flow-through select operator MUX_5289_inst
    IMA67_5290 <= type_cast_5286_wire_constant when (BITSEL_u8_u1_5284_wire(0) /=  '0') else type_cast_5288_wire_constant;
    -- logger for split-operator MUX_5299_inst flow-through 
    process(IMA68_5300) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_5299_inst:flowthrough inputs: " & " BITSEL_u8_u1_5294_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_5294_wire) & " type_cast_5296_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5296_wire_constant) & " type_cast_5298_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5298_wire_constant) & " outputs:" & " IMA68_5300= "  & Convert_SLV_To_Hex_String(IMA68_5300));
      --
    end process; 
    -- flow-through select operator MUX_5299_inst
    IMA68_5300 <= type_cast_5296_wire_constant when (BITSEL_u8_u1_5294_wire(0) /=  '0') else type_cast_5298_wire_constant;
    -- logger for split-operator MUX_5309_inst flow-through 
    process(IMA69_5310) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_5309_inst:flowthrough inputs: " & " BITSEL_u8_u1_5304_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_5304_wire) & " type_cast_5306_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5306_wire_constant) & " type_cast_5308_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5308_wire_constant) & " outputs:" & " IMA69_5310= "  & Convert_SLV_To_Hex_String(IMA69_5310));
      --
    end process; 
    -- flow-through select operator MUX_5309_inst
    IMA69_5310 <= type_cast_5306_wire_constant when (BITSEL_u8_u1_5304_wire(0) /=  '0') else type_cast_5308_wire_constant;
    -- logger for split-operator MUX_5319_inst flow-through 
    process(IMA70_5320) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_5319_inst:flowthrough inputs: " & " BITSEL_u8_u1_5314_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_5314_wire) & " type_cast_5316_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5316_wire_constant) & " type_cast_5318_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5318_wire_constant) & " outputs:" & " IMA70_5320= "  & Convert_SLV_To_Hex_String(IMA70_5320));
      --
    end process; 
    -- flow-through select operator MUX_5319_inst
    IMA70_5320 <= type_cast_5316_wire_constant when (BITSEL_u8_u1_5314_wire(0) /=  '0') else type_cast_5318_wire_constant;
    -- logger for split-operator MUX_5329_inst flow-through 
    process(IMA71_5330) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_5329_inst:flowthrough inputs: " & " BITSEL_u8_u1_5324_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_5324_wire) & " type_cast_5326_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5326_wire_constant) & " type_cast_5328_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5328_wire_constant) & " outputs:" & " IMA71_5330= "  & Convert_SLV_To_Hex_String(IMA71_5330));
      --
    end process; 
    -- flow-through select operator MUX_5329_inst
    IMA71_5330 <= type_cast_5326_wire_constant when (BITSEL_u8_u1_5324_wire(0) /=  '0') else type_cast_5328_wire_constant;
    -- logger for split-operator MUX_5339_inst flow-through 
    process(IMA72_5340) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_5339_inst:flowthrough inputs: " & " BITSEL_u8_u1_5334_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_5334_wire) & " type_cast_5336_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5336_wire_constant) & " type_cast_5338_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5338_wire_constant) & " outputs:" & " IMA72_5340= "  & Convert_SLV_To_Hex_String(IMA72_5340));
      --
    end process; 
    -- flow-through select operator MUX_5339_inst
    IMA72_5340 <= type_cast_5336_wire_constant when (BITSEL_u8_u1_5334_wire(0) /=  '0') else type_cast_5338_wire_constant;
    -- logger for split-operator MUX_5349_inst flow-through 
    process(IMA73_5350) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_5349_inst:flowthrough inputs: " & " BITSEL_u8_u1_5344_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_5344_wire) & " type_cast_5346_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5346_wire_constant) & " type_cast_5348_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5348_wire_constant) & " outputs:" & " IMA73_5350= "  & Convert_SLV_To_Hex_String(IMA73_5350));
      --
    end process; 
    -- flow-through select operator MUX_5349_inst
    IMA73_5350 <= type_cast_5346_wire_constant when (BITSEL_u8_u1_5344_wire(0) /=  '0') else type_cast_5348_wire_constant;
    -- logger for split-operator MUX_5359_inst flow-through 
    process(IMA74_5360) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_5359_inst:flowthrough inputs: " & " BITSEL_u8_u1_5354_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_5354_wire) & " type_cast_5356_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5356_wire_constant) & " type_cast_5358_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5358_wire_constant) & " outputs:" & " IMA74_5360= "  & Convert_SLV_To_Hex_String(IMA74_5360));
      --
    end process; 
    -- flow-through select operator MUX_5359_inst
    IMA74_5360 <= type_cast_5356_wire_constant when (BITSEL_u8_u1_5354_wire(0) /=  '0') else type_cast_5358_wire_constant;
    -- logger for split-operator MUX_5369_inst flow-through 
    process(IMA75_5370) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_5369_inst:flowthrough inputs: " & " BITSEL_u8_u1_5364_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_5364_wire) & " type_cast_5366_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5366_wire_constant) & " type_cast_5368_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5368_wire_constant) & " outputs:" & " IMA75_5370= "  & Convert_SLV_To_Hex_String(IMA75_5370));
      --
    end process; 
    -- flow-through select operator MUX_5369_inst
    IMA75_5370 <= type_cast_5366_wire_constant when (BITSEL_u8_u1_5364_wire(0) /=  '0') else type_cast_5368_wire_constant;
    -- logger for split-operator MUX_5379_inst flow-through 
    process(IMA76_5380) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_5379_inst:flowthrough inputs: " & " BITSEL_u8_u1_5374_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_5374_wire) & " type_cast_5376_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5376_wire_constant) & " type_cast_5378_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5378_wire_constant) & " outputs:" & " IMA76_5380= "  & Convert_SLV_To_Hex_String(IMA76_5380));
      --
    end process; 
    -- flow-through select operator MUX_5379_inst
    IMA76_5380 <= type_cast_5376_wire_constant when (BITSEL_u8_u1_5374_wire(0) /=  '0') else type_cast_5378_wire_constant;
    -- logger for split-operator MUX_5389_inst flow-through 
    process(IMA77_5390) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_5389_inst:flowthrough inputs: " & " BITSEL_u8_u1_5384_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_5384_wire) & " type_cast_5386_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5386_wire_constant) & " type_cast_5388_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5388_wire_constant) & " outputs:" & " IMA77_5390= "  & Convert_SLV_To_Hex_String(IMA77_5390));
      --
    end process; 
    -- flow-through select operator MUX_5389_inst
    IMA77_5390 <= type_cast_5386_wire_constant when (BITSEL_u8_u1_5384_wire(0) /=  '0') else type_cast_5388_wire_constant;
    -- logger for split-operator MUX_5399_inst flow-through 
    process(IMA78_5400) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_5399_inst:flowthrough inputs: " & " BITSEL_u8_u1_5394_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_5394_wire) & " type_cast_5396_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5396_wire_constant) & " type_cast_5398_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5398_wire_constant) & " outputs:" & " IMA78_5400= "  & Convert_SLV_To_Hex_String(IMA78_5400));
      --
    end process; 
    -- flow-through select operator MUX_5399_inst
    IMA78_5400 <= type_cast_5396_wire_constant when (BITSEL_u8_u1_5394_wire(0) /=  '0') else type_cast_5398_wire_constant;
    -- logger for split-operator MUX_5409_inst flow-through 
    process(IMA79_5410) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_5409_inst:flowthrough inputs: " & " BITSEL_u8_u1_5404_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_5404_wire) & " type_cast_5406_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5406_wire_constant) & " type_cast_5408_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5408_wire_constant) & " outputs:" & " IMA79_5410= "  & Convert_SLV_To_Hex_String(IMA79_5410));
      --
    end process; 
    -- flow-through select operator MUX_5409_inst
    IMA79_5410 <= type_cast_5406_wire_constant when (BITSEL_u8_u1_5404_wire(0) /=  '0') else type_cast_5408_wire_constant;
    -- logger for split-operator MUX_5419_inst flow-through 
    process(IMA80_5420) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_5419_inst:flowthrough inputs: " & " BITSEL_u8_u1_5414_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_5414_wire) & " type_cast_5416_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5416_wire_constant) & " type_cast_5418_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5418_wire_constant) & " outputs:" & " IMA80_5420= "  & Convert_SLV_To_Hex_String(IMA80_5420));
      --
    end process; 
    -- flow-through select operator MUX_5419_inst
    IMA80_5420 <= type_cast_5416_wire_constant when (BITSEL_u8_u1_5414_wire(0) /=  '0') else type_cast_5418_wire_constant;
    -- logger for split-operator MUX_5429_inst flow-through 
    process(IMA81_5430) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_5429_inst:flowthrough inputs: " & " BITSEL_u8_u1_5424_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_5424_wire) & " type_cast_5426_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5426_wire_constant) & " type_cast_5428_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5428_wire_constant) & " outputs:" & " IMA81_5430= "  & Convert_SLV_To_Hex_String(IMA81_5430));
      --
    end process; 
    -- flow-through select operator MUX_5429_inst
    IMA81_5430 <= type_cast_5426_wire_constant when (BITSEL_u8_u1_5424_wire(0) /=  '0') else type_cast_5428_wire_constant;
    -- logger for split-operator MUX_5439_inst flow-through 
    process(IMA82_5440) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_5439_inst:flowthrough inputs: " & " BITSEL_u8_u1_5434_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_5434_wire) & " type_cast_5436_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5436_wire_constant) & " type_cast_5438_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5438_wire_constant) & " outputs:" & " IMA82_5440= "  & Convert_SLV_To_Hex_String(IMA82_5440));
      --
    end process; 
    -- flow-through select operator MUX_5439_inst
    IMA82_5440 <= type_cast_5436_wire_constant when (BITSEL_u8_u1_5434_wire(0) /=  '0') else type_cast_5438_wire_constant;
    -- logger for split-operator MUX_5449_inst flow-through 
    process(IMA83_5450) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_5449_inst:flowthrough inputs: " & " BITSEL_u8_u1_5444_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_5444_wire) & " type_cast_5446_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5446_wire_constant) & " type_cast_5448_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5448_wire_constant) & " outputs:" & " IMA83_5450= "  & Convert_SLV_To_Hex_String(IMA83_5450));
      --
    end process; 
    -- flow-through select operator MUX_5449_inst
    IMA83_5450 <= type_cast_5446_wire_constant when (BITSEL_u8_u1_5444_wire(0) /=  '0') else type_cast_5448_wire_constant;
    -- logger for split-operator MUX_5459_inst flow-through 
    process(IMA84_5460) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_5459_inst:flowthrough inputs: " & " BITSEL_u8_u1_5454_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_5454_wire) & " type_cast_5456_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5456_wire_constant) & " type_cast_5458_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5458_wire_constant) & " outputs:" & " IMA84_5460= "  & Convert_SLV_To_Hex_String(IMA84_5460));
      --
    end process; 
    -- flow-through select operator MUX_5459_inst
    IMA84_5460 <= type_cast_5456_wire_constant when (BITSEL_u8_u1_5454_wire(0) /=  '0') else type_cast_5458_wire_constant;
    -- logger for split-operator MUX_5469_inst flow-through 
    process(IMA85_5470) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_5469_inst:flowthrough inputs: " & " BITSEL_u8_u1_5464_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_5464_wire) & " type_cast_5466_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5466_wire_constant) & " type_cast_5468_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5468_wire_constant) & " outputs:" & " IMA85_5470= "  & Convert_SLV_To_Hex_String(IMA85_5470));
      --
    end process; 
    -- flow-through select operator MUX_5469_inst
    IMA85_5470 <= type_cast_5466_wire_constant when (BITSEL_u8_u1_5464_wire(0) /=  '0') else type_cast_5468_wire_constant;
    -- logger for split-operator MUX_5479_inst flow-through 
    process(IMA86_5480) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_5479_inst:flowthrough inputs: " & " BITSEL_u8_u1_5474_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_5474_wire) & " type_cast_5476_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5476_wire_constant) & " type_cast_5478_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5478_wire_constant) & " outputs:" & " IMA86_5480= "  & Convert_SLV_To_Hex_String(IMA86_5480));
      --
    end process; 
    -- flow-through select operator MUX_5479_inst
    IMA86_5480 <= type_cast_5476_wire_constant when (BITSEL_u8_u1_5474_wire(0) /=  '0') else type_cast_5478_wire_constant;
    -- logger for split-operator MUX_5489_inst flow-through 
    process(IMA87_5490) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_5489_inst:flowthrough inputs: " & " BITSEL_u8_u1_5484_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_5484_wire) & " type_cast_5486_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5486_wire_constant) & " type_cast_5488_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5488_wire_constant) & " outputs:" & " IMA87_5490= "  & Convert_SLV_To_Hex_String(IMA87_5490));
      --
    end process; 
    -- flow-through select operator MUX_5489_inst
    IMA87_5490 <= type_cast_5486_wire_constant when (BITSEL_u8_u1_5484_wire(0) /=  '0') else type_cast_5488_wire_constant;
    -- logger for split-operator MUX_5499_inst flow-through 
    process(IMA88_5500) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_5499_inst:flowthrough inputs: " & " BITSEL_u8_u1_5494_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_5494_wire) & " type_cast_5496_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5496_wire_constant) & " type_cast_5498_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5498_wire_constant) & " outputs:" & " IMA88_5500= "  & Convert_SLV_To_Hex_String(IMA88_5500));
      --
    end process; 
    -- flow-through select operator MUX_5499_inst
    IMA88_5500 <= type_cast_5496_wire_constant when (BITSEL_u8_u1_5494_wire(0) /=  '0') else type_cast_5498_wire_constant;
    -- logger for split-operator MUX_5509_inst flow-through 
    process(IMA89_5510) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_5509_inst:flowthrough inputs: " & " BITSEL_u8_u1_5504_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_5504_wire) & " type_cast_5506_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5506_wire_constant) & " type_cast_5508_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5508_wire_constant) & " outputs:" & " IMA89_5510= "  & Convert_SLV_To_Hex_String(IMA89_5510));
      --
    end process; 
    -- flow-through select operator MUX_5509_inst
    IMA89_5510 <= type_cast_5506_wire_constant when (BITSEL_u8_u1_5504_wire(0) /=  '0') else type_cast_5508_wire_constant;
    -- logger for split-operator MUX_5519_inst flow-through 
    process(IMA90_5520) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_5519_inst:flowthrough inputs: " & " BITSEL_u8_u1_5514_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_5514_wire) & " type_cast_5516_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5516_wire_constant) & " type_cast_5518_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5518_wire_constant) & " outputs:" & " IMA90_5520= "  & Convert_SLV_To_Hex_String(IMA90_5520));
      --
    end process; 
    -- flow-through select operator MUX_5519_inst
    IMA90_5520 <= type_cast_5516_wire_constant when (BITSEL_u8_u1_5514_wire(0) /=  '0') else type_cast_5518_wire_constant;
    -- logger for split-operator MUX_5529_inst flow-through 
    process(IMA91_5530) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_5529_inst:flowthrough inputs: " & " BITSEL_u8_u1_5524_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_5524_wire) & " type_cast_5526_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5526_wire_constant) & " type_cast_5528_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5528_wire_constant) & " outputs:" & " IMA91_5530= "  & Convert_SLV_To_Hex_String(IMA91_5530));
      --
    end process; 
    -- flow-through select operator MUX_5529_inst
    IMA91_5530 <= type_cast_5526_wire_constant when (BITSEL_u8_u1_5524_wire(0) /=  '0') else type_cast_5528_wire_constant;
    -- logger for split-operator MUX_5539_inst flow-through 
    process(IMA92_5540) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_5539_inst:flowthrough inputs: " & " BITSEL_u8_u1_5534_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_5534_wire) & " type_cast_5536_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5536_wire_constant) & " type_cast_5538_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5538_wire_constant) & " outputs:" & " IMA92_5540= "  & Convert_SLV_To_Hex_String(IMA92_5540));
      --
    end process; 
    -- flow-through select operator MUX_5539_inst
    IMA92_5540 <= type_cast_5536_wire_constant when (BITSEL_u8_u1_5534_wire(0) /=  '0') else type_cast_5538_wire_constant;
    -- logger for split-operator MUX_5549_inst flow-through 
    process(IMA93_5550) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_5549_inst:flowthrough inputs: " & " BITSEL_u8_u1_5544_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_5544_wire) & " type_cast_5546_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5546_wire_constant) & " type_cast_5548_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5548_wire_constant) & " outputs:" & " IMA93_5550= "  & Convert_SLV_To_Hex_String(IMA93_5550));
      --
    end process; 
    -- flow-through select operator MUX_5549_inst
    IMA93_5550 <= type_cast_5546_wire_constant when (BITSEL_u8_u1_5544_wire(0) /=  '0') else type_cast_5548_wire_constant;
    -- logger for split-operator MUX_5559_inst flow-through 
    process(IMA94_5560) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_5559_inst:flowthrough inputs: " & " BITSEL_u8_u1_5554_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_5554_wire) & " type_cast_5556_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5556_wire_constant) & " type_cast_5558_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5558_wire_constant) & " outputs:" & " IMA94_5560= "  & Convert_SLV_To_Hex_String(IMA94_5560));
      --
    end process; 
    -- flow-through select operator MUX_5559_inst
    IMA94_5560 <= type_cast_5556_wire_constant when (BITSEL_u8_u1_5554_wire(0) /=  '0') else type_cast_5558_wire_constant;
    -- logger for split-operator MUX_5569_inst flow-through 
    process(IMA95_5570) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_5569_inst:flowthrough inputs: " & " BITSEL_u8_u1_5564_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_5564_wire) & " type_cast_5566_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5566_wire_constant) & " type_cast_5568_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5568_wire_constant) & " outputs:" & " IMA95_5570= "  & Convert_SLV_To_Hex_String(IMA95_5570));
      --
    end process; 
    -- flow-through select operator MUX_5569_inst
    IMA95_5570 <= type_cast_5566_wire_constant when (BITSEL_u8_u1_5564_wire(0) /=  '0') else type_cast_5568_wire_constant;
    -- logger for split-operator MUX_5579_inst flow-through 
    process(IMA96_5580) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_5579_inst:flowthrough inputs: " & " BITSEL_u8_u1_5574_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_5574_wire) & " type_cast_5576_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5576_wire_constant) & " type_cast_5578_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5578_wire_constant) & " outputs:" & " IMA96_5580= "  & Convert_SLV_To_Hex_String(IMA96_5580));
      --
    end process; 
    -- flow-through select operator MUX_5579_inst
    IMA96_5580 <= type_cast_5576_wire_constant when (BITSEL_u8_u1_5574_wire(0) /=  '0') else type_cast_5578_wire_constant;
    -- logger for split-operator MUX_5589_inst flow-through 
    process(IMA97_5590) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_5589_inst:flowthrough inputs: " & " BITSEL_u8_u1_5584_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_5584_wire) & " type_cast_5586_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5586_wire_constant) & " type_cast_5588_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5588_wire_constant) & " outputs:" & " IMA97_5590= "  & Convert_SLV_To_Hex_String(IMA97_5590));
      --
    end process; 
    -- flow-through select operator MUX_5589_inst
    IMA97_5590 <= type_cast_5586_wire_constant when (BITSEL_u8_u1_5584_wire(0) /=  '0') else type_cast_5588_wire_constant;
    -- logger for split-operator MUX_5599_inst flow-through 
    process(IMA98_5600) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_5599_inst:flowthrough inputs: " & " BITSEL_u8_u1_5594_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_5594_wire) & " type_cast_5596_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5596_wire_constant) & " type_cast_5598_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5598_wire_constant) & " outputs:" & " IMA98_5600= "  & Convert_SLV_To_Hex_String(IMA98_5600));
      --
    end process; 
    -- flow-through select operator MUX_5599_inst
    IMA98_5600 <= type_cast_5596_wire_constant when (BITSEL_u8_u1_5594_wire(0) /=  '0') else type_cast_5598_wire_constant;
    -- logger for split-operator MUX_5609_inst flow-through 
    process(IMA99_5610) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_5609_inst:flowthrough inputs: " & " BITSEL_u8_u1_5604_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_5604_wire) & " type_cast_5606_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5606_wire_constant) & " type_cast_5608_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5608_wire_constant) & " outputs:" & " IMA99_5610= "  & Convert_SLV_To_Hex_String(IMA99_5610));
      --
    end process; 
    -- flow-through select operator MUX_5609_inst
    IMA99_5610 <= type_cast_5606_wire_constant when (BITSEL_u8_u1_5604_wire(0) /=  '0') else type_cast_5608_wire_constant;
    -- logger for split-operator MUX_5619_inst flow-through 
    process(IMA100_5620) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_5619_inst:flowthrough inputs: " & " BITSEL_u8_u1_5614_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_5614_wire) & " type_cast_5616_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5616_wire_constant) & " type_cast_5618_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5618_wire_constant) & " outputs:" & " IMA100_5620= "  & Convert_SLV_To_Hex_String(IMA100_5620));
      --
    end process; 
    -- flow-through select operator MUX_5619_inst
    IMA100_5620 <= type_cast_5616_wire_constant when (BITSEL_u8_u1_5614_wire(0) /=  '0') else type_cast_5618_wire_constant;
    -- logger for split-operator MUX_5629_inst flow-through 
    process(IMA101_5630) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_5629_inst:flowthrough inputs: " & " BITSEL_u8_u1_5624_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_5624_wire) & " type_cast_5626_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5626_wire_constant) & " type_cast_5628_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5628_wire_constant) & " outputs:" & " IMA101_5630= "  & Convert_SLV_To_Hex_String(IMA101_5630));
      --
    end process; 
    -- flow-through select operator MUX_5629_inst
    IMA101_5630 <= type_cast_5626_wire_constant when (BITSEL_u8_u1_5624_wire(0) /=  '0') else type_cast_5628_wire_constant;
    -- logger for split-operator MUX_5639_inst flow-through 
    process(IMA102_5640) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_5639_inst:flowthrough inputs: " & " BITSEL_u8_u1_5634_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_5634_wire) & " type_cast_5636_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5636_wire_constant) & " type_cast_5638_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5638_wire_constant) & " outputs:" & " IMA102_5640= "  & Convert_SLV_To_Hex_String(IMA102_5640));
      --
    end process; 
    -- flow-through select operator MUX_5639_inst
    IMA102_5640 <= type_cast_5636_wire_constant when (BITSEL_u8_u1_5634_wire(0) /=  '0') else type_cast_5638_wire_constant;
    -- logger for split-operator MUX_5649_inst flow-through 
    process(IMA103_5650) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_5649_inst:flowthrough inputs: " & " BITSEL_u8_u1_5644_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_5644_wire) & " type_cast_5646_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5646_wire_constant) & " type_cast_5648_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5648_wire_constant) & " outputs:" & " IMA103_5650= "  & Convert_SLV_To_Hex_String(IMA103_5650));
      --
    end process; 
    -- flow-through select operator MUX_5649_inst
    IMA103_5650 <= type_cast_5646_wire_constant when (BITSEL_u8_u1_5644_wire(0) /=  '0') else type_cast_5648_wire_constant;
    -- logger for split-operator MUX_5659_inst flow-through 
    process(IMA104_5660) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_5659_inst:flowthrough inputs: " & " BITSEL_u8_u1_5654_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_5654_wire) & " type_cast_5656_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5656_wire_constant) & " type_cast_5658_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5658_wire_constant) & " outputs:" & " IMA104_5660= "  & Convert_SLV_To_Hex_String(IMA104_5660));
      --
    end process; 
    -- flow-through select operator MUX_5659_inst
    IMA104_5660 <= type_cast_5656_wire_constant when (BITSEL_u8_u1_5654_wire(0) /=  '0') else type_cast_5658_wire_constant;
    -- logger for split-operator MUX_5669_inst flow-through 
    process(IMA105_5670) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_5669_inst:flowthrough inputs: " & " BITSEL_u8_u1_5664_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_5664_wire) & " type_cast_5666_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5666_wire_constant) & " type_cast_5668_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5668_wire_constant) & " outputs:" & " IMA105_5670= "  & Convert_SLV_To_Hex_String(IMA105_5670));
      --
    end process; 
    -- flow-through select operator MUX_5669_inst
    IMA105_5670 <= type_cast_5666_wire_constant when (BITSEL_u8_u1_5664_wire(0) /=  '0') else type_cast_5668_wire_constant;
    -- logger for split-operator MUX_5679_inst flow-through 
    process(IMA106_5680) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_5679_inst:flowthrough inputs: " & " BITSEL_u8_u1_5674_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_5674_wire) & " type_cast_5676_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5676_wire_constant) & " type_cast_5678_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5678_wire_constant) & " outputs:" & " IMA106_5680= "  & Convert_SLV_To_Hex_String(IMA106_5680));
      --
    end process; 
    -- flow-through select operator MUX_5679_inst
    IMA106_5680 <= type_cast_5676_wire_constant when (BITSEL_u8_u1_5674_wire(0) /=  '0') else type_cast_5678_wire_constant;
    -- logger for split-operator MUX_5689_inst flow-through 
    process(IMA107_5690) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_5689_inst:flowthrough inputs: " & " BITSEL_u8_u1_5684_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_5684_wire) & " type_cast_5686_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5686_wire_constant) & " type_cast_5688_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5688_wire_constant) & " outputs:" & " IMA107_5690= "  & Convert_SLV_To_Hex_String(IMA107_5690));
      --
    end process; 
    -- flow-through select operator MUX_5689_inst
    IMA107_5690 <= type_cast_5686_wire_constant when (BITSEL_u8_u1_5684_wire(0) /=  '0') else type_cast_5688_wire_constant;
    -- logger for split-operator MUX_5699_inst flow-through 
    process(IMA108_5700) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_5699_inst:flowthrough inputs: " & " BITSEL_u8_u1_5694_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_5694_wire) & " type_cast_5696_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5696_wire_constant) & " type_cast_5698_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5698_wire_constant) & " outputs:" & " IMA108_5700= "  & Convert_SLV_To_Hex_String(IMA108_5700));
      --
    end process; 
    -- flow-through select operator MUX_5699_inst
    IMA108_5700 <= type_cast_5696_wire_constant when (BITSEL_u8_u1_5694_wire(0) /=  '0') else type_cast_5698_wire_constant;
    -- logger for split-operator MUX_5709_inst flow-through 
    process(IMA109_5710) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_5709_inst:flowthrough inputs: " & " BITSEL_u8_u1_5704_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_5704_wire) & " type_cast_5706_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5706_wire_constant) & " type_cast_5708_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5708_wire_constant) & " outputs:" & " IMA109_5710= "  & Convert_SLV_To_Hex_String(IMA109_5710));
      --
    end process; 
    -- flow-through select operator MUX_5709_inst
    IMA109_5710 <= type_cast_5706_wire_constant when (BITSEL_u8_u1_5704_wire(0) /=  '0') else type_cast_5708_wire_constant;
    -- logger for split-operator MUX_5719_inst flow-through 
    process(IMA110_5720) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_5719_inst:flowthrough inputs: " & " BITSEL_u8_u1_5714_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_5714_wire) & " type_cast_5716_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5716_wire_constant) & " type_cast_5718_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5718_wire_constant) & " outputs:" & " IMA110_5720= "  & Convert_SLV_To_Hex_String(IMA110_5720));
      --
    end process; 
    -- flow-through select operator MUX_5719_inst
    IMA110_5720 <= type_cast_5716_wire_constant when (BITSEL_u8_u1_5714_wire(0) /=  '0') else type_cast_5718_wire_constant;
    -- logger for split-operator MUX_5729_inst flow-through 
    process(IMA111_5730) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_5729_inst:flowthrough inputs: " & " BITSEL_u8_u1_5724_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_5724_wire) & " type_cast_5726_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5726_wire_constant) & " type_cast_5728_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5728_wire_constant) & " outputs:" & " IMA111_5730= "  & Convert_SLV_To_Hex_String(IMA111_5730));
      --
    end process; 
    -- flow-through select operator MUX_5729_inst
    IMA111_5730 <= type_cast_5726_wire_constant when (BITSEL_u8_u1_5724_wire(0) /=  '0') else type_cast_5728_wire_constant;
    -- logger for split-operator MUX_5739_inst flow-through 
    process(IMA112_5740) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_5739_inst:flowthrough inputs: " & " BITSEL_u8_u1_5734_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_5734_wire) & " type_cast_5736_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5736_wire_constant) & " type_cast_5738_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5738_wire_constant) & " outputs:" & " IMA112_5740= "  & Convert_SLV_To_Hex_String(IMA112_5740));
      --
    end process; 
    -- flow-through select operator MUX_5739_inst
    IMA112_5740 <= type_cast_5736_wire_constant when (BITSEL_u8_u1_5734_wire(0) /=  '0') else type_cast_5738_wire_constant;
    -- logger for split-operator MUX_5749_inst flow-through 
    process(IMA113_5750) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_5749_inst:flowthrough inputs: " & " BITSEL_u8_u1_5744_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_5744_wire) & " type_cast_5746_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5746_wire_constant) & " type_cast_5748_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5748_wire_constant) & " outputs:" & " IMA113_5750= "  & Convert_SLV_To_Hex_String(IMA113_5750));
      --
    end process; 
    -- flow-through select operator MUX_5749_inst
    IMA113_5750 <= type_cast_5746_wire_constant when (BITSEL_u8_u1_5744_wire(0) /=  '0') else type_cast_5748_wire_constant;
    -- logger for split-operator MUX_5759_inst flow-through 
    process(IMA114_5760) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_5759_inst:flowthrough inputs: " & " BITSEL_u8_u1_5754_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_5754_wire) & " type_cast_5756_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5756_wire_constant) & " type_cast_5758_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5758_wire_constant) & " outputs:" & " IMA114_5760= "  & Convert_SLV_To_Hex_String(IMA114_5760));
      --
    end process; 
    -- flow-through select operator MUX_5759_inst
    IMA114_5760 <= type_cast_5756_wire_constant when (BITSEL_u8_u1_5754_wire(0) /=  '0') else type_cast_5758_wire_constant;
    -- logger for split-operator MUX_5769_inst flow-through 
    process(IMA115_5770) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_5769_inst:flowthrough inputs: " & " BITSEL_u8_u1_5764_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_5764_wire) & " type_cast_5766_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5766_wire_constant) & " type_cast_5768_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5768_wire_constant) & " outputs:" & " IMA115_5770= "  & Convert_SLV_To_Hex_String(IMA115_5770));
      --
    end process; 
    -- flow-through select operator MUX_5769_inst
    IMA115_5770 <= type_cast_5766_wire_constant when (BITSEL_u8_u1_5764_wire(0) /=  '0') else type_cast_5768_wire_constant;
    -- logger for split-operator MUX_5779_inst flow-through 
    process(IMA116_5780) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_5779_inst:flowthrough inputs: " & " BITSEL_u8_u1_5774_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_5774_wire) & " type_cast_5776_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5776_wire_constant) & " type_cast_5778_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5778_wire_constant) & " outputs:" & " IMA116_5780= "  & Convert_SLV_To_Hex_String(IMA116_5780));
      --
    end process; 
    -- flow-through select operator MUX_5779_inst
    IMA116_5780 <= type_cast_5776_wire_constant when (BITSEL_u8_u1_5774_wire(0) /=  '0') else type_cast_5778_wire_constant;
    -- logger for split-operator MUX_5789_inst flow-through 
    process(IMA117_5790) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_5789_inst:flowthrough inputs: " & " BITSEL_u8_u1_5784_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_5784_wire) & " type_cast_5786_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5786_wire_constant) & " type_cast_5788_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5788_wire_constant) & " outputs:" & " IMA117_5790= "  & Convert_SLV_To_Hex_String(IMA117_5790));
      --
    end process; 
    -- flow-through select operator MUX_5789_inst
    IMA117_5790 <= type_cast_5786_wire_constant when (BITSEL_u8_u1_5784_wire(0) /=  '0') else type_cast_5788_wire_constant;
    -- logger for split-operator MUX_5799_inst flow-through 
    process(IMA118_5800) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_5799_inst:flowthrough inputs: " & " BITSEL_u8_u1_5794_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_5794_wire) & " type_cast_5796_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5796_wire_constant) & " type_cast_5798_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5798_wire_constant) & " outputs:" & " IMA118_5800= "  & Convert_SLV_To_Hex_String(IMA118_5800));
      --
    end process; 
    -- flow-through select operator MUX_5799_inst
    IMA118_5800 <= type_cast_5796_wire_constant when (BITSEL_u8_u1_5794_wire(0) /=  '0') else type_cast_5798_wire_constant;
    -- logger for split-operator MUX_5809_inst flow-through 
    process(IMA119_5810) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_5809_inst:flowthrough inputs: " & " BITSEL_u8_u1_5804_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_5804_wire) & " type_cast_5806_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5806_wire_constant) & " type_cast_5808_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5808_wire_constant) & " outputs:" & " IMA119_5810= "  & Convert_SLV_To_Hex_String(IMA119_5810));
      --
    end process; 
    -- flow-through select operator MUX_5809_inst
    IMA119_5810 <= type_cast_5806_wire_constant when (BITSEL_u8_u1_5804_wire(0) /=  '0') else type_cast_5808_wire_constant;
    -- logger for split-operator MUX_5819_inst flow-through 
    process(IMA120_5820) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_5819_inst:flowthrough inputs: " & " BITSEL_u8_u1_5814_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_5814_wire) & " type_cast_5816_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5816_wire_constant) & " type_cast_5818_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5818_wire_constant) & " outputs:" & " IMA120_5820= "  & Convert_SLV_To_Hex_String(IMA120_5820));
      --
    end process; 
    -- flow-through select operator MUX_5819_inst
    IMA120_5820 <= type_cast_5816_wire_constant when (BITSEL_u8_u1_5814_wire(0) /=  '0') else type_cast_5818_wire_constant;
    -- logger for split-operator MUX_5829_inst flow-through 
    process(IMA121_5830) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_5829_inst:flowthrough inputs: " & " BITSEL_u8_u1_5824_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_5824_wire) & " type_cast_5826_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5826_wire_constant) & " type_cast_5828_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5828_wire_constant) & " outputs:" & " IMA121_5830= "  & Convert_SLV_To_Hex_String(IMA121_5830));
      --
    end process; 
    -- flow-through select operator MUX_5829_inst
    IMA121_5830 <= type_cast_5826_wire_constant when (BITSEL_u8_u1_5824_wire(0) /=  '0') else type_cast_5828_wire_constant;
    -- logger for split-operator MUX_5839_inst flow-through 
    process(IMA122_5840) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_5839_inst:flowthrough inputs: " & " BITSEL_u8_u1_5834_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_5834_wire) & " type_cast_5836_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5836_wire_constant) & " type_cast_5838_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5838_wire_constant) & " outputs:" & " IMA122_5840= "  & Convert_SLV_To_Hex_String(IMA122_5840));
      --
    end process; 
    -- flow-through select operator MUX_5839_inst
    IMA122_5840 <= type_cast_5836_wire_constant when (BITSEL_u8_u1_5834_wire(0) /=  '0') else type_cast_5838_wire_constant;
    -- logger for split-operator MUX_5849_inst flow-through 
    process(IMA123_5850) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_5849_inst:flowthrough inputs: " & " BITSEL_u8_u1_5844_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_5844_wire) & " type_cast_5846_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5846_wire_constant) & " type_cast_5848_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5848_wire_constant) & " outputs:" & " IMA123_5850= "  & Convert_SLV_To_Hex_String(IMA123_5850));
      --
    end process; 
    -- flow-through select operator MUX_5849_inst
    IMA123_5850 <= type_cast_5846_wire_constant when (BITSEL_u8_u1_5844_wire(0) /=  '0') else type_cast_5848_wire_constant;
    -- logger for split-operator MUX_5859_inst flow-through 
    process(IMA124_5860) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_5859_inst:flowthrough inputs: " & " BITSEL_u8_u1_5854_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_5854_wire) & " type_cast_5856_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5856_wire_constant) & " type_cast_5858_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5858_wire_constant) & " outputs:" & " IMA124_5860= "  & Convert_SLV_To_Hex_String(IMA124_5860));
      --
    end process; 
    -- flow-through select operator MUX_5859_inst
    IMA124_5860 <= type_cast_5856_wire_constant when (BITSEL_u8_u1_5854_wire(0) /=  '0') else type_cast_5858_wire_constant;
    -- logger for split-operator MUX_5869_inst flow-through 
    process(IMA125_5870) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_5869_inst:flowthrough inputs: " & " BITSEL_u8_u1_5864_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_5864_wire) & " type_cast_5866_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5866_wire_constant) & " type_cast_5868_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5868_wire_constant) & " outputs:" & " IMA125_5870= "  & Convert_SLV_To_Hex_String(IMA125_5870));
      --
    end process; 
    -- flow-through select operator MUX_5869_inst
    IMA125_5870 <= type_cast_5866_wire_constant when (BITSEL_u8_u1_5864_wire(0) /=  '0') else type_cast_5868_wire_constant;
    -- logger for split-operator MUX_5879_inst flow-through 
    process(IMA126_5880) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_5879_inst:flowthrough inputs: " & " BITSEL_u8_u1_5874_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_5874_wire) & " type_cast_5876_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5876_wire_constant) & " type_cast_5878_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5878_wire_constant) & " outputs:" & " IMA126_5880= "  & Convert_SLV_To_Hex_String(IMA126_5880));
      --
    end process; 
    -- flow-through select operator MUX_5879_inst
    IMA126_5880 <= type_cast_5876_wire_constant when (BITSEL_u8_u1_5874_wire(0) /=  '0') else type_cast_5878_wire_constant;
    -- logger for split-operator MUX_5889_inst flow-through 
    process(IMA127_5890) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_5889_inst:flowthrough inputs: " & " BITSEL_u8_u1_5884_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_5884_wire) & " type_cast_5886_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5886_wire_constant) & " type_cast_5888_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_5888_wire_constant) & " outputs:" & " IMA127_5890= "  & Convert_SLV_To_Hex_String(IMA127_5890));
      --
    end process; 
    -- flow-through select operator MUX_5889_inst
    IMA127_5890 <= type_cast_5886_wire_constant when (BITSEL_u8_u1_5884_wire(0) /=  '0') else type_cast_5888_wire_constant;
    -- logger for split-operator MUX_5897_inst flow-through 
    process(IMB0_5898) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_5897_inst:flowthrough inputs: " & " BITSEL_u8_u1_5894_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_5894_wire) & " IMA1_4630 = "& Convert_SLV_To_Hex_String(IMA1_4630) & " IMA0_4620 = "& Convert_SLV_To_Hex_String(IMA0_4620) & " outputs:" & " IMB0_5898= "  & Convert_SLV_To_Hex_String(IMB0_5898));
      --
    end process; 
    -- flow-through select operator MUX_5897_inst
    IMB0_5898 <= IMA1_4630 when (BITSEL_u8_u1_5894_wire(0) /=  '0') else IMA0_4620;
    -- logger for split-operator MUX_5905_inst flow-through 
    process(IMB1_5906) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_5905_inst:flowthrough inputs: " & " BITSEL_u8_u1_5902_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_5902_wire) & " IMA3_4650 = "& Convert_SLV_To_Hex_String(IMA3_4650) & " IMA2_4640 = "& Convert_SLV_To_Hex_String(IMA2_4640) & " outputs:" & " IMB1_5906= "  & Convert_SLV_To_Hex_String(IMB1_5906));
      --
    end process; 
    -- flow-through select operator MUX_5905_inst
    IMB1_5906 <= IMA3_4650 when (BITSEL_u8_u1_5902_wire(0) /=  '0') else IMA2_4640;
    -- logger for split-operator MUX_5913_inst flow-through 
    process(IMB2_5914) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_5913_inst:flowthrough inputs: " & " BITSEL_u8_u1_5910_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_5910_wire) & " IMA5_4670 = "& Convert_SLV_To_Hex_String(IMA5_4670) & " IMA4_4660 = "& Convert_SLV_To_Hex_String(IMA4_4660) & " outputs:" & " IMB2_5914= "  & Convert_SLV_To_Hex_String(IMB2_5914));
      --
    end process; 
    -- flow-through select operator MUX_5913_inst
    IMB2_5914 <= IMA5_4670 when (BITSEL_u8_u1_5910_wire(0) /=  '0') else IMA4_4660;
    -- logger for split-operator MUX_5921_inst flow-through 
    process(IMB3_5922) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_5921_inst:flowthrough inputs: " & " BITSEL_u8_u1_5918_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_5918_wire) & " IMA7_4690 = "& Convert_SLV_To_Hex_String(IMA7_4690) & " IMA6_4680 = "& Convert_SLV_To_Hex_String(IMA6_4680) & " outputs:" & " IMB3_5922= "  & Convert_SLV_To_Hex_String(IMB3_5922));
      --
    end process; 
    -- flow-through select operator MUX_5921_inst
    IMB3_5922 <= IMA7_4690 when (BITSEL_u8_u1_5918_wire(0) /=  '0') else IMA6_4680;
    -- logger for split-operator MUX_5929_inst flow-through 
    process(IMB4_5930) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_5929_inst:flowthrough inputs: " & " BITSEL_u8_u1_5926_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_5926_wire) & " IMA9_4710 = "& Convert_SLV_To_Hex_String(IMA9_4710) & " IMA8_4700 = "& Convert_SLV_To_Hex_String(IMA8_4700) & " outputs:" & " IMB4_5930= "  & Convert_SLV_To_Hex_String(IMB4_5930));
      --
    end process; 
    -- flow-through select operator MUX_5929_inst
    IMB4_5930 <= IMA9_4710 when (BITSEL_u8_u1_5926_wire(0) /=  '0') else IMA8_4700;
    -- logger for split-operator MUX_5937_inst flow-through 
    process(IMB5_5938) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_5937_inst:flowthrough inputs: " & " BITSEL_u8_u1_5934_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_5934_wire) & " IMA11_4730 = "& Convert_SLV_To_Hex_String(IMA11_4730) & " IMA10_4720 = "& Convert_SLV_To_Hex_String(IMA10_4720) & " outputs:" & " IMB5_5938= "  & Convert_SLV_To_Hex_String(IMB5_5938));
      --
    end process; 
    -- flow-through select operator MUX_5937_inst
    IMB5_5938 <= IMA11_4730 when (BITSEL_u8_u1_5934_wire(0) /=  '0') else IMA10_4720;
    -- logger for split-operator MUX_5945_inst flow-through 
    process(IMB6_5946) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_5945_inst:flowthrough inputs: " & " BITSEL_u8_u1_5942_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_5942_wire) & " IMA13_4750 = "& Convert_SLV_To_Hex_String(IMA13_4750) & " IMA12_4740 = "& Convert_SLV_To_Hex_String(IMA12_4740) & " outputs:" & " IMB6_5946= "  & Convert_SLV_To_Hex_String(IMB6_5946));
      --
    end process; 
    -- flow-through select operator MUX_5945_inst
    IMB6_5946 <= IMA13_4750 when (BITSEL_u8_u1_5942_wire(0) /=  '0') else IMA12_4740;
    -- logger for split-operator MUX_5953_inst flow-through 
    process(IMB7_5954) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_5953_inst:flowthrough inputs: " & " BITSEL_u8_u1_5950_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_5950_wire) & " IMA15_4770 = "& Convert_SLV_To_Hex_String(IMA15_4770) & " IMA14_4760 = "& Convert_SLV_To_Hex_String(IMA14_4760) & " outputs:" & " IMB7_5954= "  & Convert_SLV_To_Hex_String(IMB7_5954));
      --
    end process; 
    -- flow-through select operator MUX_5953_inst
    IMB7_5954 <= IMA15_4770 when (BITSEL_u8_u1_5950_wire(0) /=  '0') else IMA14_4760;
    -- logger for split-operator MUX_5961_inst flow-through 
    process(IMB8_5962) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_5961_inst:flowthrough inputs: " & " BITSEL_u8_u1_5958_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_5958_wire) & " IMA17_4790 = "& Convert_SLV_To_Hex_String(IMA17_4790) & " IMA16_4780 = "& Convert_SLV_To_Hex_String(IMA16_4780) & " outputs:" & " IMB8_5962= "  & Convert_SLV_To_Hex_String(IMB8_5962));
      --
    end process; 
    -- flow-through select operator MUX_5961_inst
    IMB8_5962 <= IMA17_4790 when (BITSEL_u8_u1_5958_wire(0) /=  '0') else IMA16_4780;
    -- logger for split-operator MUX_5969_inst flow-through 
    process(IMB9_5970) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_5969_inst:flowthrough inputs: " & " BITSEL_u8_u1_5966_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_5966_wire) & " IMA19_4810 = "& Convert_SLV_To_Hex_String(IMA19_4810) & " IMA18_4800 = "& Convert_SLV_To_Hex_String(IMA18_4800) & " outputs:" & " IMB9_5970= "  & Convert_SLV_To_Hex_String(IMB9_5970));
      --
    end process; 
    -- flow-through select operator MUX_5969_inst
    IMB9_5970 <= IMA19_4810 when (BITSEL_u8_u1_5966_wire(0) /=  '0') else IMA18_4800;
    -- logger for split-operator MUX_5977_inst flow-through 
    process(IMB10_5978) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_5977_inst:flowthrough inputs: " & " BITSEL_u8_u1_5974_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_5974_wire) & " IMA21_4830 = "& Convert_SLV_To_Hex_String(IMA21_4830) & " IMA20_4820 = "& Convert_SLV_To_Hex_String(IMA20_4820) & " outputs:" & " IMB10_5978= "  & Convert_SLV_To_Hex_String(IMB10_5978));
      --
    end process; 
    -- flow-through select operator MUX_5977_inst
    IMB10_5978 <= IMA21_4830 when (BITSEL_u8_u1_5974_wire(0) /=  '0') else IMA20_4820;
    -- logger for split-operator MUX_5985_inst flow-through 
    process(IMB11_5986) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_5985_inst:flowthrough inputs: " & " BITSEL_u8_u1_5982_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_5982_wire) & " IMA23_4850 = "& Convert_SLV_To_Hex_String(IMA23_4850) & " IMA22_4840 = "& Convert_SLV_To_Hex_String(IMA22_4840) & " outputs:" & " IMB11_5986= "  & Convert_SLV_To_Hex_String(IMB11_5986));
      --
    end process; 
    -- flow-through select operator MUX_5985_inst
    IMB11_5986 <= IMA23_4850 when (BITSEL_u8_u1_5982_wire(0) /=  '0') else IMA22_4840;
    -- logger for split-operator MUX_5993_inst flow-through 
    process(IMB12_5994) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_5993_inst:flowthrough inputs: " & " BITSEL_u8_u1_5990_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_5990_wire) & " IMA25_4870 = "& Convert_SLV_To_Hex_String(IMA25_4870) & " IMA24_4860 = "& Convert_SLV_To_Hex_String(IMA24_4860) & " outputs:" & " IMB12_5994= "  & Convert_SLV_To_Hex_String(IMB12_5994));
      --
    end process; 
    -- flow-through select operator MUX_5993_inst
    IMB12_5994 <= IMA25_4870 when (BITSEL_u8_u1_5990_wire(0) /=  '0') else IMA24_4860;
    -- logger for split-operator MUX_6001_inst flow-through 
    process(IMB13_6002) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6001_inst:flowthrough inputs: " & " BITSEL_u8_u1_5998_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_5998_wire) & " IMA27_4890 = "& Convert_SLV_To_Hex_String(IMA27_4890) & " IMA26_4880 = "& Convert_SLV_To_Hex_String(IMA26_4880) & " outputs:" & " IMB13_6002= "  & Convert_SLV_To_Hex_String(IMB13_6002));
      --
    end process; 
    -- flow-through select operator MUX_6001_inst
    IMB13_6002 <= IMA27_4890 when (BITSEL_u8_u1_5998_wire(0) /=  '0') else IMA26_4880;
    -- logger for split-operator MUX_6009_inst flow-through 
    process(IMB14_6010) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6009_inst:flowthrough inputs: " & " BITSEL_u8_u1_6006_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6006_wire) & " IMA29_4910 = "& Convert_SLV_To_Hex_String(IMA29_4910) & " IMA28_4900 = "& Convert_SLV_To_Hex_String(IMA28_4900) & " outputs:" & " IMB14_6010= "  & Convert_SLV_To_Hex_String(IMB14_6010));
      --
    end process; 
    -- flow-through select operator MUX_6009_inst
    IMB14_6010 <= IMA29_4910 when (BITSEL_u8_u1_6006_wire(0) /=  '0') else IMA28_4900;
    -- logger for split-operator MUX_6017_inst flow-through 
    process(IMB15_6018) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6017_inst:flowthrough inputs: " & " BITSEL_u8_u1_6014_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6014_wire) & " IMA31_4930 = "& Convert_SLV_To_Hex_String(IMA31_4930) & " IMA30_4920 = "& Convert_SLV_To_Hex_String(IMA30_4920) & " outputs:" & " IMB15_6018= "  & Convert_SLV_To_Hex_String(IMB15_6018));
      --
    end process; 
    -- flow-through select operator MUX_6017_inst
    IMB15_6018 <= IMA31_4930 when (BITSEL_u8_u1_6014_wire(0) /=  '0') else IMA30_4920;
    -- logger for split-operator MUX_6025_inst flow-through 
    process(IMB16_6026) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6025_inst:flowthrough inputs: " & " BITSEL_u8_u1_6022_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6022_wire) & " IMA33_4950 = "& Convert_SLV_To_Hex_String(IMA33_4950) & " IMA32_4940 = "& Convert_SLV_To_Hex_String(IMA32_4940) & " outputs:" & " IMB16_6026= "  & Convert_SLV_To_Hex_String(IMB16_6026));
      --
    end process; 
    -- flow-through select operator MUX_6025_inst
    IMB16_6026 <= IMA33_4950 when (BITSEL_u8_u1_6022_wire(0) /=  '0') else IMA32_4940;
    -- logger for split-operator MUX_6033_inst flow-through 
    process(IMB17_6034) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6033_inst:flowthrough inputs: " & " BITSEL_u8_u1_6030_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6030_wire) & " IMA35_4970 = "& Convert_SLV_To_Hex_String(IMA35_4970) & " IMA34_4960 = "& Convert_SLV_To_Hex_String(IMA34_4960) & " outputs:" & " IMB17_6034= "  & Convert_SLV_To_Hex_String(IMB17_6034));
      --
    end process; 
    -- flow-through select operator MUX_6033_inst
    IMB17_6034 <= IMA35_4970 when (BITSEL_u8_u1_6030_wire(0) /=  '0') else IMA34_4960;
    -- logger for split-operator MUX_6041_inst flow-through 
    process(IMB18_6042) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6041_inst:flowthrough inputs: " & " BITSEL_u8_u1_6038_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6038_wire) & " IMA37_4990 = "& Convert_SLV_To_Hex_String(IMA37_4990) & " IMA36_4980 = "& Convert_SLV_To_Hex_String(IMA36_4980) & " outputs:" & " IMB18_6042= "  & Convert_SLV_To_Hex_String(IMB18_6042));
      --
    end process; 
    -- flow-through select operator MUX_6041_inst
    IMB18_6042 <= IMA37_4990 when (BITSEL_u8_u1_6038_wire(0) /=  '0') else IMA36_4980;
    -- logger for split-operator MUX_6049_inst flow-through 
    process(IMB19_6050) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6049_inst:flowthrough inputs: " & " BITSEL_u8_u1_6046_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6046_wire) & " IMA39_5010 = "& Convert_SLV_To_Hex_String(IMA39_5010) & " IMA38_5000 = "& Convert_SLV_To_Hex_String(IMA38_5000) & " outputs:" & " IMB19_6050= "  & Convert_SLV_To_Hex_String(IMB19_6050));
      --
    end process; 
    -- flow-through select operator MUX_6049_inst
    IMB19_6050 <= IMA39_5010 when (BITSEL_u8_u1_6046_wire(0) /=  '0') else IMA38_5000;
    -- logger for split-operator MUX_6057_inst flow-through 
    process(IMB20_6058) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6057_inst:flowthrough inputs: " & " BITSEL_u8_u1_6054_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6054_wire) & " IMA41_5030 = "& Convert_SLV_To_Hex_String(IMA41_5030) & " IMA40_5020 = "& Convert_SLV_To_Hex_String(IMA40_5020) & " outputs:" & " IMB20_6058= "  & Convert_SLV_To_Hex_String(IMB20_6058));
      --
    end process; 
    -- flow-through select operator MUX_6057_inst
    IMB20_6058 <= IMA41_5030 when (BITSEL_u8_u1_6054_wire(0) /=  '0') else IMA40_5020;
    -- logger for split-operator MUX_6065_inst flow-through 
    process(IMB21_6066) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6065_inst:flowthrough inputs: " & " BITSEL_u8_u1_6062_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6062_wire) & " IMA43_5050 = "& Convert_SLV_To_Hex_String(IMA43_5050) & " IMA42_5040 = "& Convert_SLV_To_Hex_String(IMA42_5040) & " outputs:" & " IMB21_6066= "  & Convert_SLV_To_Hex_String(IMB21_6066));
      --
    end process; 
    -- flow-through select operator MUX_6065_inst
    IMB21_6066 <= IMA43_5050 when (BITSEL_u8_u1_6062_wire(0) /=  '0') else IMA42_5040;
    -- logger for split-operator MUX_6073_inst flow-through 
    process(IMB22_6074) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6073_inst:flowthrough inputs: " & " BITSEL_u8_u1_6070_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6070_wire) & " IMA45_5070 = "& Convert_SLV_To_Hex_String(IMA45_5070) & " IMA44_5060 = "& Convert_SLV_To_Hex_String(IMA44_5060) & " outputs:" & " IMB22_6074= "  & Convert_SLV_To_Hex_String(IMB22_6074));
      --
    end process; 
    -- flow-through select operator MUX_6073_inst
    IMB22_6074 <= IMA45_5070 when (BITSEL_u8_u1_6070_wire(0) /=  '0') else IMA44_5060;
    -- logger for split-operator MUX_6081_inst flow-through 
    process(IMB23_6082) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6081_inst:flowthrough inputs: " & " BITSEL_u8_u1_6078_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6078_wire) & " IMA47_5090 = "& Convert_SLV_To_Hex_String(IMA47_5090) & " IMA46_5080 = "& Convert_SLV_To_Hex_String(IMA46_5080) & " outputs:" & " IMB23_6082= "  & Convert_SLV_To_Hex_String(IMB23_6082));
      --
    end process; 
    -- flow-through select operator MUX_6081_inst
    IMB23_6082 <= IMA47_5090 when (BITSEL_u8_u1_6078_wire(0) /=  '0') else IMA46_5080;
    -- logger for split-operator MUX_6089_inst flow-through 
    process(IMB24_6090) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6089_inst:flowthrough inputs: " & " BITSEL_u8_u1_6086_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6086_wire) & " IMA49_5110 = "& Convert_SLV_To_Hex_String(IMA49_5110) & " IMA48_5100 = "& Convert_SLV_To_Hex_String(IMA48_5100) & " outputs:" & " IMB24_6090= "  & Convert_SLV_To_Hex_String(IMB24_6090));
      --
    end process; 
    -- flow-through select operator MUX_6089_inst
    IMB24_6090 <= IMA49_5110 when (BITSEL_u8_u1_6086_wire(0) /=  '0') else IMA48_5100;
    -- logger for split-operator MUX_6097_inst flow-through 
    process(IMB25_6098) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6097_inst:flowthrough inputs: " & " BITSEL_u8_u1_6094_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6094_wire) & " IMA51_5130 = "& Convert_SLV_To_Hex_String(IMA51_5130) & " IMA50_5120 = "& Convert_SLV_To_Hex_String(IMA50_5120) & " outputs:" & " IMB25_6098= "  & Convert_SLV_To_Hex_String(IMB25_6098));
      --
    end process; 
    -- flow-through select operator MUX_6097_inst
    IMB25_6098 <= IMA51_5130 when (BITSEL_u8_u1_6094_wire(0) /=  '0') else IMA50_5120;
    -- logger for split-operator MUX_6105_inst flow-through 
    process(IMB26_6106) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6105_inst:flowthrough inputs: " & " BITSEL_u8_u1_6102_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6102_wire) & " IMA53_5150 = "& Convert_SLV_To_Hex_String(IMA53_5150) & " IMA52_5140 = "& Convert_SLV_To_Hex_String(IMA52_5140) & " outputs:" & " IMB26_6106= "  & Convert_SLV_To_Hex_String(IMB26_6106));
      --
    end process; 
    -- flow-through select operator MUX_6105_inst
    IMB26_6106 <= IMA53_5150 when (BITSEL_u8_u1_6102_wire(0) /=  '0') else IMA52_5140;
    -- logger for split-operator MUX_6113_inst flow-through 
    process(IMB27_6114) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6113_inst:flowthrough inputs: " & " BITSEL_u8_u1_6110_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6110_wire) & " IMA55_5170 = "& Convert_SLV_To_Hex_String(IMA55_5170) & " IMA54_5160 = "& Convert_SLV_To_Hex_String(IMA54_5160) & " outputs:" & " IMB27_6114= "  & Convert_SLV_To_Hex_String(IMB27_6114));
      --
    end process; 
    -- flow-through select operator MUX_6113_inst
    IMB27_6114 <= IMA55_5170 when (BITSEL_u8_u1_6110_wire(0) /=  '0') else IMA54_5160;
    -- logger for split-operator MUX_6121_inst flow-through 
    process(IMB28_6122) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6121_inst:flowthrough inputs: " & " BITSEL_u8_u1_6118_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6118_wire) & " IMA57_5190 = "& Convert_SLV_To_Hex_String(IMA57_5190) & " IMA56_5180 = "& Convert_SLV_To_Hex_String(IMA56_5180) & " outputs:" & " IMB28_6122= "  & Convert_SLV_To_Hex_String(IMB28_6122));
      --
    end process; 
    -- flow-through select operator MUX_6121_inst
    IMB28_6122 <= IMA57_5190 when (BITSEL_u8_u1_6118_wire(0) /=  '0') else IMA56_5180;
    -- logger for split-operator MUX_6129_inst flow-through 
    process(IMB29_6130) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6129_inst:flowthrough inputs: " & " BITSEL_u8_u1_6126_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6126_wire) & " IMA59_5210 = "& Convert_SLV_To_Hex_String(IMA59_5210) & " IMA58_5200 = "& Convert_SLV_To_Hex_String(IMA58_5200) & " outputs:" & " IMB29_6130= "  & Convert_SLV_To_Hex_String(IMB29_6130));
      --
    end process; 
    -- flow-through select operator MUX_6129_inst
    IMB29_6130 <= IMA59_5210 when (BITSEL_u8_u1_6126_wire(0) /=  '0') else IMA58_5200;
    -- logger for split-operator MUX_6137_inst flow-through 
    process(IMB30_6138) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6137_inst:flowthrough inputs: " & " BITSEL_u8_u1_6134_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6134_wire) & " IMA61_5230 = "& Convert_SLV_To_Hex_String(IMA61_5230) & " IMA60_5220 = "& Convert_SLV_To_Hex_String(IMA60_5220) & " outputs:" & " IMB30_6138= "  & Convert_SLV_To_Hex_String(IMB30_6138));
      --
    end process; 
    -- flow-through select operator MUX_6137_inst
    IMB30_6138 <= IMA61_5230 when (BITSEL_u8_u1_6134_wire(0) /=  '0') else IMA60_5220;
    -- logger for split-operator MUX_6145_inst flow-through 
    process(IMB31_6146) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6145_inst:flowthrough inputs: " & " BITSEL_u8_u1_6142_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6142_wire) & " IMA63_5250 = "& Convert_SLV_To_Hex_String(IMA63_5250) & " IMA62_5240 = "& Convert_SLV_To_Hex_String(IMA62_5240) & " outputs:" & " IMB31_6146= "  & Convert_SLV_To_Hex_String(IMB31_6146));
      --
    end process; 
    -- flow-through select operator MUX_6145_inst
    IMB31_6146 <= IMA63_5250 when (BITSEL_u8_u1_6142_wire(0) /=  '0') else IMA62_5240;
    -- logger for split-operator MUX_6153_inst flow-through 
    process(IMB32_6154) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6153_inst:flowthrough inputs: " & " BITSEL_u8_u1_6150_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6150_wire) & " IMA65_5270 = "& Convert_SLV_To_Hex_String(IMA65_5270) & " IMA64_5260 = "& Convert_SLV_To_Hex_String(IMA64_5260) & " outputs:" & " IMB32_6154= "  & Convert_SLV_To_Hex_String(IMB32_6154));
      --
    end process; 
    -- flow-through select operator MUX_6153_inst
    IMB32_6154 <= IMA65_5270 when (BITSEL_u8_u1_6150_wire(0) /=  '0') else IMA64_5260;
    -- logger for split-operator MUX_6161_inst flow-through 
    process(IMB33_6162) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6161_inst:flowthrough inputs: " & " BITSEL_u8_u1_6158_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6158_wire) & " IMA67_5290 = "& Convert_SLV_To_Hex_String(IMA67_5290) & " IMA66_5280 = "& Convert_SLV_To_Hex_String(IMA66_5280) & " outputs:" & " IMB33_6162= "  & Convert_SLV_To_Hex_String(IMB33_6162));
      --
    end process; 
    -- flow-through select operator MUX_6161_inst
    IMB33_6162 <= IMA67_5290 when (BITSEL_u8_u1_6158_wire(0) /=  '0') else IMA66_5280;
    -- logger for split-operator MUX_6169_inst flow-through 
    process(IMB34_6170) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6169_inst:flowthrough inputs: " & " BITSEL_u8_u1_6166_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6166_wire) & " IMA69_5310 = "& Convert_SLV_To_Hex_String(IMA69_5310) & " IMA68_5300 = "& Convert_SLV_To_Hex_String(IMA68_5300) & " outputs:" & " IMB34_6170= "  & Convert_SLV_To_Hex_String(IMB34_6170));
      --
    end process; 
    -- flow-through select operator MUX_6169_inst
    IMB34_6170 <= IMA69_5310 when (BITSEL_u8_u1_6166_wire(0) /=  '0') else IMA68_5300;
    -- logger for split-operator MUX_6177_inst flow-through 
    process(IMB35_6178) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6177_inst:flowthrough inputs: " & " BITSEL_u8_u1_6174_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6174_wire) & " IMA71_5330 = "& Convert_SLV_To_Hex_String(IMA71_5330) & " IMA70_5320 = "& Convert_SLV_To_Hex_String(IMA70_5320) & " outputs:" & " IMB35_6178= "  & Convert_SLV_To_Hex_String(IMB35_6178));
      --
    end process; 
    -- flow-through select operator MUX_6177_inst
    IMB35_6178 <= IMA71_5330 when (BITSEL_u8_u1_6174_wire(0) /=  '0') else IMA70_5320;
    -- logger for split-operator MUX_6185_inst flow-through 
    process(IMB36_6186) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6185_inst:flowthrough inputs: " & " BITSEL_u8_u1_6182_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6182_wire) & " IMA73_5350 = "& Convert_SLV_To_Hex_String(IMA73_5350) & " IMA72_5340 = "& Convert_SLV_To_Hex_String(IMA72_5340) & " outputs:" & " IMB36_6186= "  & Convert_SLV_To_Hex_String(IMB36_6186));
      --
    end process; 
    -- flow-through select operator MUX_6185_inst
    IMB36_6186 <= IMA73_5350 when (BITSEL_u8_u1_6182_wire(0) /=  '0') else IMA72_5340;
    -- logger for split-operator MUX_6193_inst flow-through 
    process(IMB37_6194) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6193_inst:flowthrough inputs: " & " BITSEL_u8_u1_6190_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6190_wire) & " IMA75_5370 = "& Convert_SLV_To_Hex_String(IMA75_5370) & " IMA74_5360 = "& Convert_SLV_To_Hex_String(IMA74_5360) & " outputs:" & " IMB37_6194= "  & Convert_SLV_To_Hex_String(IMB37_6194));
      --
    end process; 
    -- flow-through select operator MUX_6193_inst
    IMB37_6194 <= IMA75_5370 when (BITSEL_u8_u1_6190_wire(0) /=  '0') else IMA74_5360;
    -- logger for split-operator MUX_6201_inst flow-through 
    process(IMB38_6202) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6201_inst:flowthrough inputs: " & " BITSEL_u8_u1_6198_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6198_wire) & " IMA77_5390 = "& Convert_SLV_To_Hex_String(IMA77_5390) & " IMA76_5380 = "& Convert_SLV_To_Hex_String(IMA76_5380) & " outputs:" & " IMB38_6202= "  & Convert_SLV_To_Hex_String(IMB38_6202));
      --
    end process; 
    -- flow-through select operator MUX_6201_inst
    IMB38_6202 <= IMA77_5390 when (BITSEL_u8_u1_6198_wire(0) /=  '0') else IMA76_5380;
    -- logger for split-operator MUX_6209_inst flow-through 
    process(IMB39_6210) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6209_inst:flowthrough inputs: " & " BITSEL_u8_u1_6206_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6206_wire) & " IMA79_5410 = "& Convert_SLV_To_Hex_String(IMA79_5410) & " IMA78_5400 = "& Convert_SLV_To_Hex_String(IMA78_5400) & " outputs:" & " IMB39_6210= "  & Convert_SLV_To_Hex_String(IMB39_6210));
      --
    end process; 
    -- flow-through select operator MUX_6209_inst
    IMB39_6210 <= IMA79_5410 when (BITSEL_u8_u1_6206_wire(0) /=  '0') else IMA78_5400;
    -- logger for split-operator MUX_6217_inst flow-through 
    process(IMB40_6218) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6217_inst:flowthrough inputs: " & " BITSEL_u8_u1_6214_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6214_wire) & " IMA81_5430 = "& Convert_SLV_To_Hex_String(IMA81_5430) & " IMA80_5420 = "& Convert_SLV_To_Hex_String(IMA80_5420) & " outputs:" & " IMB40_6218= "  & Convert_SLV_To_Hex_String(IMB40_6218));
      --
    end process; 
    -- flow-through select operator MUX_6217_inst
    IMB40_6218 <= IMA81_5430 when (BITSEL_u8_u1_6214_wire(0) /=  '0') else IMA80_5420;
    -- logger for split-operator MUX_6225_inst flow-through 
    process(IMB41_6226) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6225_inst:flowthrough inputs: " & " BITSEL_u8_u1_6222_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6222_wire) & " IMA83_5450 = "& Convert_SLV_To_Hex_String(IMA83_5450) & " IMA82_5440 = "& Convert_SLV_To_Hex_String(IMA82_5440) & " outputs:" & " IMB41_6226= "  & Convert_SLV_To_Hex_String(IMB41_6226));
      --
    end process; 
    -- flow-through select operator MUX_6225_inst
    IMB41_6226 <= IMA83_5450 when (BITSEL_u8_u1_6222_wire(0) /=  '0') else IMA82_5440;
    -- logger for split-operator MUX_6233_inst flow-through 
    process(IMB42_6234) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6233_inst:flowthrough inputs: " & " BITSEL_u8_u1_6230_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6230_wire) & " IMA85_5470 = "& Convert_SLV_To_Hex_String(IMA85_5470) & " IMA84_5460 = "& Convert_SLV_To_Hex_String(IMA84_5460) & " outputs:" & " IMB42_6234= "  & Convert_SLV_To_Hex_String(IMB42_6234));
      --
    end process; 
    -- flow-through select operator MUX_6233_inst
    IMB42_6234 <= IMA85_5470 when (BITSEL_u8_u1_6230_wire(0) /=  '0') else IMA84_5460;
    -- logger for split-operator MUX_6241_inst flow-through 
    process(IMB43_6242) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6241_inst:flowthrough inputs: " & " BITSEL_u8_u1_6238_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6238_wire) & " IMA87_5490 = "& Convert_SLV_To_Hex_String(IMA87_5490) & " IMA86_5480 = "& Convert_SLV_To_Hex_String(IMA86_5480) & " outputs:" & " IMB43_6242= "  & Convert_SLV_To_Hex_String(IMB43_6242));
      --
    end process; 
    -- flow-through select operator MUX_6241_inst
    IMB43_6242 <= IMA87_5490 when (BITSEL_u8_u1_6238_wire(0) /=  '0') else IMA86_5480;
    -- logger for split-operator MUX_6249_inst flow-through 
    process(IMB44_6250) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6249_inst:flowthrough inputs: " & " BITSEL_u8_u1_6246_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6246_wire) & " IMA89_5510 = "& Convert_SLV_To_Hex_String(IMA89_5510) & " IMA88_5500 = "& Convert_SLV_To_Hex_String(IMA88_5500) & " outputs:" & " IMB44_6250= "  & Convert_SLV_To_Hex_String(IMB44_6250));
      --
    end process; 
    -- flow-through select operator MUX_6249_inst
    IMB44_6250 <= IMA89_5510 when (BITSEL_u8_u1_6246_wire(0) /=  '0') else IMA88_5500;
    -- logger for split-operator MUX_6257_inst flow-through 
    process(IMB45_6258) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6257_inst:flowthrough inputs: " & " BITSEL_u8_u1_6254_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6254_wire) & " IMA91_5530 = "& Convert_SLV_To_Hex_String(IMA91_5530) & " IMA90_5520 = "& Convert_SLV_To_Hex_String(IMA90_5520) & " outputs:" & " IMB45_6258= "  & Convert_SLV_To_Hex_String(IMB45_6258));
      --
    end process; 
    -- flow-through select operator MUX_6257_inst
    IMB45_6258 <= IMA91_5530 when (BITSEL_u8_u1_6254_wire(0) /=  '0') else IMA90_5520;
    -- logger for split-operator MUX_6265_inst flow-through 
    process(IMB46_6266) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6265_inst:flowthrough inputs: " & " BITSEL_u8_u1_6262_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6262_wire) & " IMA93_5550 = "& Convert_SLV_To_Hex_String(IMA93_5550) & " IMA92_5540 = "& Convert_SLV_To_Hex_String(IMA92_5540) & " outputs:" & " IMB46_6266= "  & Convert_SLV_To_Hex_String(IMB46_6266));
      --
    end process; 
    -- flow-through select operator MUX_6265_inst
    IMB46_6266 <= IMA93_5550 when (BITSEL_u8_u1_6262_wire(0) /=  '0') else IMA92_5540;
    -- logger for split-operator MUX_6273_inst flow-through 
    process(IMB47_6274) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6273_inst:flowthrough inputs: " & " BITSEL_u8_u1_6270_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6270_wire) & " IMA95_5570 = "& Convert_SLV_To_Hex_String(IMA95_5570) & " IMA94_5560 = "& Convert_SLV_To_Hex_String(IMA94_5560) & " outputs:" & " IMB47_6274= "  & Convert_SLV_To_Hex_String(IMB47_6274));
      --
    end process; 
    -- flow-through select operator MUX_6273_inst
    IMB47_6274 <= IMA95_5570 when (BITSEL_u8_u1_6270_wire(0) /=  '0') else IMA94_5560;
    -- logger for split-operator MUX_6281_inst flow-through 
    process(IMB48_6282) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6281_inst:flowthrough inputs: " & " BITSEL_u8_u1_6278_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6278_wire) & " IMA97_5590 = "& Convert_SLV_To_Hex_String(IMA97_5590) & " IMA96_5580 = "& Convert_SLV_To_Hex_String(IMA96_5580) & " outputs:" & " IMB48_6282= "  & Convert_SLV_To_Hex_String(IMB48_6282));
      --
    end process; 
    -- flow-through select operator MUX_6281_inst
    IMB48_6282 <= IMA97_5590 when (BITSEL_u8_u1_6278_wire(0) /=  '0') else IMA96_5580;
    -- logger for split-operator MUX_6289_inst flow-through 
    process(IMB49_6290) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6289_inst:flowthrough inputs: " & " BITSEL_u8_u1_6286_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6286_wire) & " IMA99_5610 = "& Convert_SLV_To_Hex_String(IMA99_5610) & " IMA98_5600 = "& Convert_SLV_To_Hex_String(IMA98_5600) & " outputs:" & " IMB49_6290= "  & Convert_SLV_To_Hex_String(IMB49_6290));
      --
    end process; 
    -- flow-through select operator MUX_6289_inst
    IMB49_6290 <= IMA99_5610 when (BITSEL_u8_u1_6286_wire(0) /=  '0') else IMA98_5600;
    -- logger for split-operator MUX_6297_inst flow-through 
    process(IMB50_6298) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6297_inst:flowthrough inputs: " & " BITSEL_u8_u1_6294_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6294_wire) & " IMA101_5630 = "& Convert_SLV_To_Hex_String(IMA101_5630) & " IMA100_5620 = "& Convert_SLV_To_Hex_String(IMA100_5620) & " outputs:" & " IMB50_6298= "  & Convert_SLV_To_Hex_String(IMB50_6298));
      --
    end process; 
    -- flow-through select operator MUX_6297_inst
    IMB50_6298 <= IMA101_5630 when (BITSEL_u8_u1_6294_wire(0) /=  '0') else IMA100_5620;
    -- logger for split-operator MUX_6305_inst flow-through 
    process(IMB51_6306) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6305_inst:flowthrough inputs: " & " BITSEL_u8_u1_6302_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6302_wire) & " IMA103_5650 = "& Convert_SLV_To_Hex_String(IMA103_5650) & " IMA102_5640 = "& Convert_SLV_To_Hex_String(IMA102_5640) & " outputs:" & " IMB51_6306= "  & Convert_SLV_To_Hex_String(IMB51_6306));
      --
    end process; 
    -- flow-through select operator MUX_6305_inst
    IMB51_6306 <= IMA103_5650 when (BITSEL_u8_u1_6302_wire(0) /=  '0') else IMA102_5640;
    -- logger for split-operator MUX_6313_inst flow-through 
    process(IMB52_6314) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6313_inst:flowthrough inputs: " & " BITSEL_u8_u1_6310_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6310_wire) & " IMA105_5670 = "& Convert_SLV_To_Hex_String(IMA105_5670) & " IMA104_5660 = "& Convert_SLV_To_Hex_String(IMA104_5660) & " outputs:" & " IMB52_6314= "  & Convert_SLV_To_Hex_String(IMB52_6314));
      --
    end process; 
    -- flow-through select operator MUX_6313_inst
    IMB52_6314 <= IMA105_5670 when (BITSEL_u8_u1_6310_wire(0) /=  '0') else IMA104_5660;
    -- logger for split-operator MUX_6321_inst flow-through 
    process(IMB53_6322) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6321_inst:flowthrough inputs: " & " BITSEL_u8_u1_6318_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6318_wire) & " IMA107_5690 = "& Convert_SLV_To_Hex_String(IMA107_5690) & " IMA106_5680 = "& Convert_SLV_To_Hex_String(IMA106_5680) & " outputs:" & " IMB53_6322= "  & Convert_SLV_To_Hex_String(IMB53_6322));
      --
    end process; 
    -- flow-through select operator MUX_6321_inst
    IMB53_6322 <= IMA107_5690 when (BITSEL_u8_u1_6318_wire(0) /=  '0') else IMA106_5680;
    -- logger for split-operator MUX_6329_inst flow-through 
    process(IMB54_6330) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6329_inst:flowthrough inputs: " & " BITSEL_u8_u1_6326_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6326_wire) & " IMA109_5710 = "& Convert_SLV_To_Hex_String(IMA109_5710) & " IMA108_5700 = "& Convert_SLV_To_Hex_String(IMA108_5700) & " outputs:" & " IMB54_6330= "  & Convert_SLV_To_Hex_String(IMB54_6330));
      --
    end process; 
    -- flow-through select operator MUX_6329_inst
    IMB54_6330 <= IMA109_5710 when (BITSEL_u8_u1_6326_wire(0) /=  '0') else IMA108_5700;
    -- logger for split-operator MUX_6337_inst flow-through 
    process(IMB55_6338) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6337_inst:flowthrough inputs: " & " BITSEL_u8_u1_6334_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6334_wire) & " IMA111_5730 = "& Convert_SLV_To_Hex_String(IMA111_5730) & " IMA110_5720 = "& Convert_SLV_To_Hex_String(IMA110_5720) & " outputs:" & " IMB55_6338= "  & Convert_SLV_To_Hex_String(IMB55_6338));
      --
    end process; 
    -- flow-through select operator MUX_6337_inst
    IMB55_6338 <= IMA111_5730 when (BITSEL_u8_u1_6334_wire(0) /=  '0') else IMA110_5720;
    -- logger for split-operator MUX_6345_inst flow-through 
    process(IMB56_6346) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6345_inst:flowthrough inputs: " & " BITSEL_u8_u1_6342_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6342_wire) & " IMA113_5750 = "& Convert_SLV_To_Hex_String(IMA113_5750) & " IMA112_5740 = "& Convert_SLV_To_Hex_String(IMA112_5740) & " outputs:" & " IMB56_6346= "  & Convert_SLV_To_Hex_String(IMB56_6346));
      --
    end process; 
    -- flow-through select operator MUX_6345_inst
    IMB56_6346 <= IMA113_5750 when (BITSEL_u8_u1_6342_wire(0) /=  '0') else IMA112_5740;
    -- logger for split-operator MUX_6353_inst flow-through 
    process(IMB57_6354) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6353_inst:flowthrough inputs: " & " BITSEL_u8_u1_6350_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6350_wire) & " IMA115_5770 = "& Convert_SLV_To_Hex_String(IMA115_5770) & " IMA114_5760 = "& Convert_SLV_To_Hex_String(IMA114_5760) & " outputs:" & " IMB57_6354= "  & Convert_SLV_To_Hex_String(IMB57_6354));
      --
    end process; 
    -- flow-through select operator MUX_6353_inst
    IMB57_6354 <= IMA115_5770 when (BITSEL_u8_u1_6350_wire(0) /=  '0') else IMA114_5760;
    -- logger for split-operator MUX_6361_inst flow-through 
    process(IMB58_6362) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6361_inst:flowthrough inputs: " & " BITSEL_u8_u1_6358_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6358_wire) & " IMA117_5790 = "& Convert_SLV_To_Hex_String(IMA117_5790) & " IMA116_5780 = "& Convert_SLV_To_Hex_String(IMA116_5780) & " outputs:" & " IMB58_6362= "  & Convert_SLV_To_Hex_String(IMB58_6362));
      --
    end process; 
    -- flow-through select operator MUX_6361_inst
    IMB58_6362 <= IMA117_5790 when (BITSEL_u8_u1_6358_wire(0) /=  '0') else IMA116_5780;
    -- logger for split-operator MUX_6369_inst flow-through 
    process(IMB59_6370) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6369_inst:flowthrough inputs: " & " BITSEL_u8_u1_6366_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6366_wire) & " IMA119_5810 = "& Convert_SLV_To_Hex_String(IMA119_5810) & " IMA118_5800 = "& Convert_SLV_To_Hex_String(IMA118_5800) & " outputs:" & " IMB59_6370= "  & Convert_SLV_To_Hex_String(IMB59_6370));
      --
    end process; 
    -- flow-through select operator MUX_6369_inst
    IMB59_6370 <= IMA119_5810 when (BITSEL_u8_u1_6366_wire(0) /=  '0') else IMA118_5800;
    -- logger for split-operator MUX_6377_inst flow-through 
    process(IMB60_6378) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6377_inst:flowthrough inputs: " & " BITSEL_u8_u1_6374_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6374_wire) & " IMA121_5830 = "& Convert_SLV_To_Hex_String(IMA121_5830) & " IMA120_5820 = "& Convert_SLV_To_Hex_String(IMA120_5820) & " outputs:" & " IMB60_6378= "  & Convert_SLV_To_Hex_String(IMB60_6378));
      --
    end process; 
    -- flow-through select operator MUX_6377_inst
    IMB60_6378 <= IMA121_5830 when (BITSEL_u8_u1_6374_wire(0) /=  '0') else IMA120_5820;
    -- logger for split-operator MUX_6385_inst flow-through 
    process(IMB61_6386) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6385_inst:flowthrough inputs: " & " BITSEL_u8_u1_6382_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6382_wire) & " IMA123_5850 = "& Convert_SLV_To_Hex_String(IMA123_5850) & " IMA122_5840 = "& Convert_SLV_To_Hex_String(IMA122_5840) & " outputs:" & " IMB61_6386= "  & Convert_SLV_To_Hex_String(IMB61_6386));
      --
    end process; 
    -- flow-through select operator MUX_6385_inst
    IMB61_6386 <= IMA123_5850 when (BITSEL_u8_u1_6382_wire(0) /=  '0') else IMA122_5840;
    -- logger for split-operator MUX_6393_inst flow-through 
    process(IMB62_6394) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6393_inst:flowthrough inputs: " & " BITSEL_u8_u1_6390_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6390_wire) & " IMA125_5870 = "& Convert_SLV_To_Hex_String(IMA125_5870) & " IMA124_5860 = "& Convert_SLV_To_Hex_String(IMA124_5860) & " outputs:" & " IMB62_6394= "  & Convert_SLV_To_Hex_String(IMB62_6394));
      --
    end process; 
    -- flow-through select operator MUX_6393_inst
    IMB62_6394 <= IMA125_5870 when (BITSEL_u8_u1_6390_wire(0) /=  '0') else IMA124_5860;
    -- logger for split-operator MUX_6401_inst flow-through 
    process(IMB63_6402) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6401_inst:flowthrough inputs: " & " BITSEL_u8_u1_6398_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6398_wire) & " IMA127_5890 = "& Convert_SLV_To_Hex_String(IMA127_5890) & " IMA126_5880 = "& Convert_SLV_To_Hex_String(IMA126_5880) & " outputs:" & " IMB63_6402= "  & Convert_SLV_To_Hex_String(IMB63_6402));
      --
    end process; 
    -- flow-through select operator MUX_6401_inst
    IMB63_6402 <= IMA127_5890 when (BITSEL_u8_u1_6398_wire(0) /=  '0') else IMA126_5880;
    -- logger for split-operator MUX_6409_inst flow-through 
    process(IMC0_6410) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6409_inst:flowthrough inputs: " & " BITSEL_u8_u1_6406_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6406_wire) & " IMB1_5906 = "& Convert_SLV_To_Hex_String(IMB1_5906) & " IMB0_5898 = "& Convert_SLV_To_Hex_String(IMB0_5898) & " outputs:" & " IMC0_6410= "  & Convert_SLV_To_Hex_String(IMC0_6410));
      --
    end process; 
    -- flow-through select operator MUX_6409_inst
    IMC0_6410 <= IMB1_5906 when (BITSEL_u8_u1_6406_wire(0) /=  '0') else IMB0_5898;
    -- logger for split-operator MUX_6417_inst flow-through 
    process(IMC1_6418) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6417_inst:flowthrough inputs: " & " BITSEL_u8_u1_6414_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6414_wire) & " IMB3_5922 = "& Convert_SLV_To_Hex_String(IMB3_5922) & " IMB2_5914 = "& Convert_SLV_To_Hex_String(IMB2_5914) & " outputs:" & " IMC1_6418= "  & Convert_SLV_To_Hex_String(IMC1_6418));
      --
    end process; 
    -- flow-through select operator MUX_6417_inst
    IMC1_6418 <= IMB3_5922 when (BITSEL_u8_u1_6414_wire(0) /=  '0') else IMB2_5914;
    -- logger for split-operator MUX_6425_inst flow-through 
    process(IMC2_6426) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6425_inst:flowthrough inputs: " & " BITSEL_u8_u1_6422_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6422_wire) & " IMB5_5938 = "& Convert_SLV_To_Hex_String(IMB5_5938) & " IMB4_5930 = "& Convert_SLV_To_Hex_String(IMB4_5930) & " outputs:" & " IMC2_6426= "  & Convert_SLV_To_Hex_String(IMC2_6426));
      --
    end process; 
    -- flow-through select operator MUX_6425_inst
    IMC2_6426 <= IMB5_5938 when (BITSEL_u8_u1_6422_wire(0) /=  '0') else IMB4_5930;
    -- logger for split-operator MUX_6433_inst flow-through 
    process(IMC3_6434) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6433_inst:flowthrough inputs: " & " BITSEL_u8_u1_6430_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6430_wire) & " IMB7_5954 = "& Convert_SLV_To_Hex_String(IMB7_5954) & " IMB6_5946 = "& Convert_SLV_To_Hex_String(IMB6_5946) & " outputs:" & " IMC3_6434= "  & Convert_SLV_To_Hex_String(IMC3_6434));
      --
    end process; 
    -- flow-through select operator MUX_6433_inst
    IMC3_6434 <= IMB7_5954 when (BITSEL_u8_u1_6430_wire(0) /=  '0') else IMB6_5946;
    -- logger for split-operator MUX_6441_inst flow-through 
    process(IMC4_6442) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6441_inst:flowthrough inputs: " & " BITSEL_u8_u1_6438_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6438_wire) & " IMB9_5970 = "& Convert_SLV_To_Hex_String(IMB9_5970) & " IMB8_5962 = "& Convert_SLV_To_Hex_String(IMB8_5962) & " outputs:" & " IMC4_6442= "  & Convert_SLV_To_Hex_String(IMC4_6442));
      --
    end process; 
    -- flow-through select operator MUX_6441_inst
    IMC4_6442 <= IMB9_5970 when (BITSEL_u8_u1_6438_wire(0) /=  '0') else IMB8_5962;
    -- logger for split-operator MUX_6449_inst flow-through 
    process(IMC5_6450) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6449_inst:flowthrough inputs: " & " BITSEL_u8_u1_6446_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6446_wire) & " IMB11_5986 = "& Convert_SLV_To_Hex_String(IMB11_5986) & " IMB10_5978 = "& Convert_SLV_To_Hex_String(IMB10_5978) & " outputs:" & " IMC5_6450= "  & Convert_SLV_To_Hex_String(IMC5_6450));
      --
    end process; 
    -- flow-through select operator MUX_6449_inst
    IMC5_6450 <= IMB11_5986 when (BITSEL_u8_u1_6446_wire(0) /=  '0') else IMB10_5978;
    -- logger for split-operator MUX_6457_inst flow-through 
    process(IMC6_6458) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6457_inst:flowthrough inputs: " & " BITSEL_u8_u1_6454_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6454_wire) & " IMB13_6002 = "& Convert_SLV_To_Hex_String(IMB13_6002) & " IMB12_5994 = "& Convert_SLV_To_Hex_String(IMB12_5994) & " outputs:" & " IMC6_6458= "  & Convert_SLV_To_Hex_String(IMC6_6458));
      --
    end process; 
    -- flow-through select operator MUX_6457_inst
    IMC6_6458 <= IMB13_6002 when (BITSEL_u8_u1_6454_wire(0) /=  '0') else IMB12_5994;
    -- logger for split-operator MUX_6465_inst flow-through 
    process(IMC7_6466) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6465_inst:flowthrough inputs: " & " BITSEL_u8_u1_6462_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6462_wire) & " IMB15_6018 = "& Convert_SLV_To_Hex_String(IMB15_6018) & " IMB14_6010 = "& Convert_SLV_To_Hex_String(IMB14_6010) & " outputs:" & " IMC7_6466= "  & Convert_SLV_To_Hex_String(IMC7_6466));
      --
    end process; 
    -- flow-through select operator MUX_6465_inst
    IMC7_6466 <= IMB15_6018 when (BITSEL_u8_u1_6462_wire(0) /=  '0') else IMB14_6010;
    -- logger for split-operator MUX_6473_inst flow-through 
    process(IMC8_6474) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6473_inst:flowthrough inputs: " & " BITSEL_u8_u1_6470_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6470_wire) & " IMB17_6034 = "& Convert_SLV_To_Hex_String(IMB17_6034) & " IMB16_6026 = "& Convert_SLV_To_Hex_String(IMB16_6026) & " outputs:" & " IMC8_6474= "  & Convert_SLV_To_Hex_String(IMC8_6474));
      --
    end process; 
    -- flow-through select operator MUX_6473_inst
    IMC8_6474 <= IMB17_6034 when (BITSEL_u8_u1_6470_wire(0) /=  '0') else IMB16_6026;
    -- logger for split-operator MUX_6481_inst flow-through 
    process(IMC9_6482) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6481_inst:flowthrough inputs: " & " BITSEL_u8_u1_6478_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6478_wire) & " IMB19_6050 = "& Convert_SLV_To_Hex_String(IMB19_6050) & " IMB18_6042 = "& Convert_SLV_To_Hex_String(IMB18_6042) & " outputs:" & " IMC9_6482= "  & Convert_SLV_To_Hex_String(IMC9_6482));
      --
    end process; 
    -- flow-through select operator MUX_6481_inst
    IMC9_6482 <= IMB19_6050 when (BITSEL_u8_u1_6478_wire(0) /=  '0') else IMB18_6042;
    -- logger for split-operator MUX_6489_inst flow-through 
    process(IMC10_6490) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6489_inst:flowthrough inputs: " & " BITSEL_u8_u1_6486_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6486_wire) & " IMB21_6066 = "& Convert_SLV_To_Hex_String(IMB21_6066) & " IMB20_6058 = "& Convert_SLV_To_Hex_String(IMB20_6058) & " outputs:" & " IMC10_6490= "  & Convert_SLV_To_Hex_String(IMC10_6490));
      --
    end process; 
    -- flow-through select operator MUX_6489_inst
    IMC10_6490 <= IMB21_6066 when (BITSEL_u8_u1_6486_wire(0) /=  '0') else IMB20_6058;
    -- logger for split-operator MUX_6497_inst flow-through 
    process(IMC11_6498) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6497_inst:flowthrough inputs: " & " BITSEL_u8_u1_6494_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6494_wire) & " IMB23_6082 = "& Convert_SLV_To_Hex_String(IMB23_6082) & " IMB22_6074 = "& Convert_SLV_To_Hex_String(IMB22_6074) & " outputs:" & " IMC11_6498= "  & Convert_SLV_To_Hex_String(IMC11_6498));
      --
    end process; 
    -- flow-through select operator MUX_6497_inst
    IMC11_6498 <= IMB23_6082 when (BITSEL_u8_u1_6494_wire(0) /=  '0') else IMB22_6074;
    -- logger for split-operator MUX_6505_inst flow-through 
    process(IMC12_6506) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6505_inst:flowthrough inputs: " & " BITSEL_u8_u1_6502_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6502_wire) & " IMB25_6098 = "& Convert_SLV_To_Hex_String(IMB25_6098) & " IMB24_6090 = "& Convert_SLV_To_Hex_String(IMB24_6090) & " outputs:" & " IMC12_6506= "  & Convert_SLV_To_Hex_String(IMC12_6506));
      --
    end process; 
    -- flow-through select operator MUX_6505_inst
    IMC12_6506 <= IMB25_6098 when (BITSEL_u8_u1_6502_wire(0) /=  '0') else IMB24_6090;
    -- logger for split-operator MUX_6513_inst flow-through 
    process(IMC13_6514) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6513_inst:flowthrough inputs: " & " BITSEL_u8_u1_6510_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6510_wire) & " IMB27_6114 = "& Convert_SLV_To_Hex_String(IMB27_6114) & " IMB26_6106 = "& Convert_SLV_To_Hex_String(IMB26_6106) & " outputs:" & " IMC13_6514= "  & Convert_SLV_To_Hex_String(IMC13_6514));
      --
    end process; 
    -- flow-through select operator MUX_6513_inst
    IMC13_6514 <= IMB27_6114 when (BITSEL_u8_u1_6510_wire(0) /=  '0') else IMB26_6106;
    -- logger for split-operator MUX_6521_inst flow-through 
    process(IMC14_6522) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6521_inst:flowthrough inputs: " & " BITSEL_u8_u1_6518_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6518_wire) & " IMB29_6130 = "& Convert_SLV_To_Hex_String(IMB29_6130) & " IMB28_6122 = "& Convert_SLV_To_Hex_String(IMB28_6122) & " outputs:" & " IMC14_6522= "  & Convert_SLV_To_Hex_String(IMC14_6522));
      --
    end process; 
    -- flow-through select operator MUX_6521_inst
    IMC14_6522 <= IMB29_6130 when (BITSEL_u8_u1_6518_wire(0) /=  '0') else IMB28_6122;
    -- logger for split-operator MUX_6529_inst flow-through 
    process(IMC15_6530) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6529_inst:flowthrough inputs: " & " BITSEL_u8_u1_6526_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6526_wire) & " IMB31_6146 = "& Convert_SLV_To_Hex_String(IMB31_6146) & " IMB30_6138 = "& Convert_SLV_To_Hex_String(IMB30_6138) & " outputs:" & " IMC15_6530= "  & Convert_SLV_To_Hex_String(IMC15_6530));
      --
    end process; 
    -- flow-through select operator MUX_6529_inst
    IMC15_6530 <= IMB31_6146 when (BITSEL_u8_u1_6526_wire(0) /=  '0') else IMB30_6138;
    -- logger for split-operator MUX_6537_inst flow-through 
    process(IMC16_6538) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6537_inst:flowthrough inputs: " & " BITSEL_u8_u1_6534_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6534_wire) & " IMB33_6162 = "& Convert_SLV_To_Hex_String(IMB33_6162) & " IMB32_6154 = "& Convert_SLV_To_Hex_String(IMB32_6154) & " outputs:" & " IMC16_6538= "  & Convert_SLV_To_Hex_String(IMC16_6538));
      --
    end process; 
    -- flow-through select operator MUX_6537_inst
    IMC16_6538 <= IMB33_6162 when (BITSEL_u8_u1_6534_wire(0) /=  '0') else IMB32_6154;
    -- logger for split-operator MUX_6545_inst flow-through 
    process(IMC17_6546) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6545_inst:flowthrough inputs: " & " BITSEL_u8_u1_6542_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6542_wire) & " IMB35_6178 = "& Convert_SLV_To_Hex_String(IMB35_6178) & " IMB34_6170 = "& Convert_SLV_To_Hex_String(IMB34_6170) & " outputs:" & " IMC17_6546= "  & Convert_SLV_To_Hex_String(IMC17_6546));
      --
    end process; 
    -- flow-through select operator MUX_6545_inst
    IMC17_6546 <= IMB35_6178 when (BITSEL_u8_u1_6542_wire(0) /=  '0') else IMB34_6170;
    -- logger for split-operator MUX_6553_inst flow-through 
    process(IMC18_6554) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6553_inst:flowthrough inputs: " & " BITSEL_u8_u1_6550_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6550_wire) & " IMB37_6194 = "& Convert_SLV_To_Hex_String(IMB37_6194) & " IMB36_6186 = "& Convert_SLV_To_Hex_String(IMB36_6186) & " outputs:" & " IMC18_6554= "  & Convert_SLV_To_Hex_String(IMC18_6554));
      --
    end process; 
    -- flow-through select operator MUX_6553_inst
    IMC18_6554 <= IMB37_6194 when (BITSEL_u8_u1_6550_wire(0) /=  '0') else IMB36_6186;
    -- logger for split-operator MUX_6561_inst flow-through 
    process(IMC19_6562) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6561_inst:flowthrough inputs: " & " BITSEL_u8_u1_6558_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6558_wire) & " IMB39_6210 = "& Convert_SLV_To_Hex_String(IMB39_6210) & " IMB38_6202 = "& Convert_SLV_To_Hex_String(IMB38_6202) & " outputs:" & " IMC19_6562= "  & Convert_SLV_To_Hex_String(IMC19_6562));
      --
    end process; 
    -- flow-through select operator MUX_6561_inst
    IMC19_6562 <= IMB39_6210 when (BITSEL_u8_u1_6558_wire(0) /=  '0') else IMB38_6202;
    -- logger for split-operator MUX_6569_inst flow-through 
    process(IMC20_6570) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6569_inst:flowthrough inputs: " & " BITSEL_u8_u1_6566_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6566_wire) & " IMB41_6226 = "& Convert_SLV_To_Hex_String(IMB41_6226) & " IMB40_6218 = "& Convert_SLV_To_Hex_String(IMB40_6218) & " outputs:" & " IMC20_6570= "  & Convert_SLV_To_Hex_String(IMC20_6570));
      --
    end process; 
    -- flow-through select operator MUX_6569_inst
    IMC20_6570 <= IMB41_6226 when (BITSEL_u8_u1_6566_wire(0) /=  '0') else IMB40_6218;
    -- logger for split-operator MUX_6577_inst flow-through 
    process(IMC21_6578) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6577_inst:flowthrough inputs: " & " BITSEL_u8_u1_6574_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6574_wire) & " IMB43_6242 = "& Convert_SLV_To_Hex_String(IMB43_6242) & " IMB42_6234 = "& Convert_SLV_To_Hex_String(IMB42_6234) & " outputs:" & " IMC21_6578= "  & Convert_SLV_To_Hex_String(IMC21_6578));
      --
    end process; 
    -- flow-through select operator MUX_6577_inst
    IMC21_6578 <= IMB43_6242 when (BITSEL_u8_u1_6574_wire(0) /=  '0') else IMB42_6234;
    -- logger for split-operator MUX_6585_inst flow-through 
    process(IMC22_6586) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6585_inst:flowthrough inputs: " & " BITSEL_u8_u1_6582_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6582_wire) & " IMB45_6258 = "& Convert_SLV_To_Hex_String(IMB45_6258) & " IMB44_6250 = "& Convert_SLV_To_Hex_String(IMB44_6250) & " outputs:" & " IMC22_6586= "  & Convert_SLV_To_Hex_String(IMC22_6586));
      --
    end process; 
    -- flow-through select operator MUX_6585_inst
    IMC22_6586 <= IMB45_6258 when (BITSEL_u8_u1_6582_wire(0) /=  '0') else IMB44_6250;
    -- logger for split-operator MUX_6593_inst flow-through 
    process(IMC23_6594) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6593_inst:flowthrough inputs: " & " BITSEL_u8_u1_6590_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6590_wire) & " IMB47_6274 = "& Convert_SLV_To_Hex_String(IMB47_6274) & " IMB46_6266 = "& Convert_SLV_To_Hex_String(IMB46_6266) & " outputs:" & " IMC23_6594= "  & Convert_SLV_To_Hex_String(IMC23_6594));
      --
    end process; 
    -- flow-through select operator MUX_6593_inst
    IMC23_6594 <= IMB47_6274 when (BITSEL_u8_u1_6590_wire(0) /=  '0') else IMB46_6266;
    -- logger for split-operator MUX_6601_inst flow-through 
    process(IMC24_6602) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6601_inst:flowthrough inputs: " & " BITSEL_u8_u1_6598_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6598_wire) & " IMB49_6290 = "& Convert_SLV_To_Hex_String(IMB49_6290) & " IMB48_6282 = "& Convert_SLV_To_Hex_String(IMB48_6282) & " outputs:" & " IMC24_6602= "  & Convert_SLV_To_Hex_String(IMC24_6602));
      --
    end process; 
    -- flow-through select operator MUX_6601_inst
    IMC24_6602 <= IMB49_6290 when (BITSEL_u8_u1_6598_wire(0) /=  '0') else IMB48_6282;
    -- logger for split-operator MUX_6609_inst flow-through 
    process(IMC25_6610) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6609_inst:flowthrough inputs: " & " BITSEL_u8_u1_6606_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6606_wire) & " IMB51_6306 = "& Convert_SLV_To_Hex_String(IMB51_6306) & " IMB50_6298 = "& Convert_SLV_To_Hex_String(IMB50_6298) & " outputs:" & " IMC25_6610= "  & Convert_SLV_To_Hex_String(IMC25_6610));
      --
    end process; 
    -- flow-through select operator MUX_6609_inst
    IMC25_6610 <= IMB51_6306 when (BITSEL_u8_u1_6606_wire(0) /=  '0') else IMB50_6298;
    -- logger for split-operator MUX_6617_inst flow-through 
    process(IMC26_6618) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6617_inst:flowthrough inputs: " & " BITSEL_u8_u1_6614_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6614_wire) & " IMB53_6322 = "& Convert_SLV_To_Hex_String(IMB53_6322) & " IMB52_6314 = "& Convert_SLV_To_Hex_String(IMB52_6314) & " outputs:" & " IMC26_6618= "  & Convert_SLV_To_Hex_String(IMC26_6618));
      --
    end process; 
    -- flow-through select operator MUX_6617_inst
    IMC26_6618 <= IMB53_6322 when (BITSEL_u8_u1_6614_wire(0) /=  '0') else IMB52_6314;
    -- logger for split-operator MUX_6625_inst flow-through 
    process(IMC27_6626) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6625_inst:flowthrough inputs: " & " BITSEL_u8_u1_6622_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6622_wire) & " IMB55_6338 = "& Convert_SLV_To_Hex_String(IMB55_6338) & " IMB54_6330 = "& Convert_SLV_To_Hex_String(IMB54_6330) & " outputs:" & " IMC27_6626= "  & Convert_SLV_To_Hex_String(IMC27_6626));
      --
    end process; 
    -- flow-through select operator MUX_6625_inst
    IMC27_6626 <= IMB55_6338 when (BITSEL_u8_u1_6622_wire(0) /=  '0') else IMB54_6330;
    -- logger for split-operator MUX_6633_inst flow-through 
    process(IMC28_6634) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6633_inst:flowthrough inputs: " & " BITSEL_u8_u1_6630_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6630_wire) & " IMB57_6354 = "& Convert_SLV_To_Hex_String(IMB57_6354) & " IMB56_6346 = "& Convert_SLV_To_Hex_String(IMB56_6346) & " outputs:" & " IMC28_6634= "  & Convert_SLV_To_Hex_String(IMC28_6634));
      --
    end process; 
    -- flow-through select operator MUX_6633_inst
    IMC28_6634 <= IMB57_6354 when (BITSEL_u8_u1_6630_wire(0) /=  '0') else IMB56_6346;
    -- logger for split-operator MUX_6641_inst flow-through 
    process(IMC29_6642) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6641_inst:flowthrough inputs: " & " BITSEL_u8_u1_6638_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6638_wire) & " IMB59_6370 = "& Convert_SLV_To_Hex_String(IMB59_6370) & " IMB58_6362 = "& Convert_SLV_To_Hex_String(IMB58_6362) & " outputs:" & " IMC29_6642= "  & Convert_SLV_To_Hex_String(IMC29_6642));
      --
    end process; 
    -- flow-through select operator MUX_6641_inst
    IMC29_6642 <= IMB59_6370 when (BITSEL_u8_u1_6638_wire(0) /=  '0') else IMB58_6362;
    -- logger for split-operator MUX_6649_inst flow-through 
    process(IMC30_6650) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6649_inst:flowthrough inputs: " & " BITSEL_u8_u1_6646_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6646_wire) & " IMB61_6386 = "& Convert_SLV_To_Hex_String(IMB61_6386) & " IMB60_6378 = "& Convert_SLV_To_Hex_String(IMB60_6378) & " outputs:" & " IMC30_6650= "  & Convert_SLV_To_Hex_String(IMC30_6650));
      --
    end process; 
    -- flow-through select operator MUX_6649_inst
    IMC30_6650 <= IMB61_6386 when (BITSEL_u8_u1_6646_wire(0) /=  '0') else IMB60_6378;
    -- logger for split-operator MUX_6657_inst flow-through 
    process(IMC31_6658) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6657_inst:flowthrough inputs: " & " BITSEL_u8_u1_6654_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6654_wire) & " IMB63_6402 = "& Convert_SLV_To_Hex_String(IMB63_6402) & " IMB62_6394 = "& Convert_SLV_To_Hex_String(IMB62_6394) & " outputs:" & " IMC31_6658= "  & Convert_SLV_To_Hex_String(IMC31_6658));
      --
    end process; 
    -- flow-through select operator MUX_6657_inst
    IMC31_6658 <= IMB63_6402 when (BITSEL_u8_u1_6654_wire(0) /=  '0') else IMB62_6394;
    -- logger for split-operator MUX_6665_inst flow-through 
    process(IMD0_6666) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6665_inst:flowthrough inputs: " & " BITSEL_u8_u1_6662_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6662_wire) & " IMC1_6418 = "& Convert_SLV_To_Hex_String(IMC1_6418) & " IMC0_6410 = "& Convert_SLV_To_Hex_String(IMC0_6410) & " outputs:" & " IMD0_6666= "  & Convert_SLV_To_Hex_String(IMD0_6666));
      --
    end process; 
    -- flow-through select operator MUX_6665_inst
    IMD0_6666 <= IMC1_6418 when (BITSEL_u8_u1_6662_wire(0) /=  '0') else IMC0_6410;
    -- logger for split-operator MUX_6673_inst flow-through 
    process(IMD1_6674) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6673_inst:flowthrough inputs: " & " BITSEL_u8_u1_6670_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6670_wire) & " IMC3_6434 = "& Convert_SLV_To_Hex_String(IMC3_6434) & " IMC2_6426 = "& Convert_SLV_To_Hex_String(IMC2_6426) & " outputs:" & " IMD1_6674= "  & Convert_SLV_To_Hex_String(IMD1_6674));
      --
    end process; 
    -- flow-through select operator MUX_6673_inst
    IMD1_6674 <= IMC3_6434 when (BITSEL_u8_u1_6670_wire(0) /=  '0') else IMC2_6426;
    -- logger for split-operator MUX_6681_inst flow-through 
    process(IMD2_6682) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6681_inst:flowthrough inputs: " & " BITSEL_u8_u1_6678_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6678_wire) & " IMC5_6450 = "& Convert_SLV_To_Hex_String(IMC5_6450) & " IMC4_6442 = "& Convert_SLV_To_Hex_String(IMC4_6442) & " outputs:" & " IMD2_6682= "  & Convert_SLV_To_Hex_String(IMD2_6682));
      --
    end process; 
    -- flow-through select operator MUX_6681_inst
    IMD2_6682 <= IMC5_6450 when (BITSEL_u8_u1_6678_wire(0) /=  '0') else IMC4_6442;
    -- logger for split-operator MUX_6689_inst flow-through 
    process(IMD3_6690) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6689_inst:flowthrough inputs: " & " BITSEL_u8_u1_6686_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6686_wire) & " IMC7_6466 = "& Convert_SLV_To_Hex_String(IMC7_6466) & " IMC6_6458 = "& Convert_SLV_To_Hex_String(IMC6_6458) & " outputs:" & " IMD3_6690= "  & Convert_SLV_To_Hex_String(IMD3_6690));
      --
    end process; 
    -- flow-through select operator MUX_6689_inst
    IMD3_6690 <= IMC7_6466 when (BITSEL_u8_u1_6686_wire(0) /=  '0') else IMC6_6458;
    -- logger for split-operator MUX_6697_inst flow-through 
    process(IMD4_6698) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6697_inst:flowthrough inputs: " & " BITSEL_u8_u1_6694_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6694_wire) & " IMC9_6482 = "& Convert_SLV_To_Hex_String(IMC9_6482) & " IMC8_6474 = "& Convert_SLV_To_Hex_String(IMC8_6474) & " outputs:" & " IMD4_6698= "  & Convert_SLV_To_Hex_String(IMD4_6698));
      --
    end process; 
    -- flow-through select operator MUX_6697_inst
    IMD4_6698 <= IMC9_6482 when (BITSEL_u8_u1_6694_wire(0) /=  '0') else IMC8_6474;
    -- logger for split-operator MUX_6705_inst flow-through 
    process(IMD5_6706) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6705_inst:flowthrough inputs: " & " BITSEL_u8_u1_6702_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6702_wire) & " IMC11_6498 = "& Convert_SLV_To_Hex_String(IMC11_6498) & " IMC10_6490 = "& Convert_SLV_To_Hex_String(IMC10_6490) & " outputs:" & " IMD5_6706= "  & Convert_SLV_To_Hex_String(IMD5_6706));
      --
    end process; 
    -- flow-through select operator MUX_6705_inst
    IMD5_6706 <= IMC11_6498 when (BITSEL_u8_u1_6702_wire(0) /=  '0') else IMC10_6490;
    -- logger for split-operator MUX_6713_inst flow-through 
    process(IMD6_6714) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6713_inst:flowthrough inputs: " & " BITSEL_u8_u1_6710_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6710_wire) & " IMC13_6514 = "& Convert_SLV_To_Hex_String(IMC13_6514) & " IMC12_6506 = "& Convert_SLV_To_Hex_String(IMC12_6506) & " outputs:" & " IMD6_6714= "  & Convert_SLV_To_Hex_String(IMD6_6714));
      --
    end process; 
    -- flow-through select operator MUX_6713_inst
    IMD6_6714 <= IMC13_6514 when (BITSEL_u8_u1_6710_wire(0) /=  '0') else IMC12_6506;
    -- logger for split-operator MUX_6721_inst flow-through 
    process(IMD7_6722) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6721_inst:flowthrough inputs: " & " BITSEL_u8_u1_6718_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6718_wire) & " IMC15_6530 = "& Convert_SLV_To_Hex_String(IMC15_6530) & " IMC14_6522 = "& Convert_SLV_To_Hex_String(IMC14_6522) & " outputs:" & " IMD7_6722= "  & Convert_SLV_To_Hex_String(IMD7_6722));
      --
    end process; 
    -- flow-through select operator MUX_6721_inst
    IMD7_6722 <= IMC15_6530 when (BITSEL_u8_u1_6718_wire(0) /=  '0') else IMC14_6522;
    -- logger for split-operator MUX_6729_inst flow-through 
    process(IMD8_6730) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6729_inst:flowthrough inputs: " & " BITSEL_u8_u1_6726_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6726_wire) & " IMC17_6546 = "& Convert_SLV_To_Hex_String(IMC17_6546) & " IMC16_6538 = "& Convert_SLV_To_Hex_String(IMC16_6538) & " outputs:" & " IMD8_6730= "  & Convert_SLV_To_Hex_String(IMD8_6730));
      --
    end process; 
    -- flow-through select operator MUX_6729_inst
    IMD8_6730 <= IMC17_6546 when (BITSEL_u8_u1_6726_wire(0) /=  '0') else IMC16_6538;
    -- logger for split-operator MUX_6737_inst flow-through 
    process(IMD9_6738) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6737_inst:flowthrough inputs: " & " BITSEL_u8_u1_6734_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6734_wire) & " IMC19_6562 = "& Convert_SLV_To_Hex_String(IMC19_6562) & " IMC18_6554 = "& Convert_SLV_To_Hex_String(IMC18_6554) & " outputs:" & " IMD9_6738= "  & Convert_SLV_To_Hex_String(IMD9_6738));
      --
    end process; 
    -- flow-through select operator MUX_6737_inst
    IMD9_6738 <= IMC19_6562 when (BITSEL_u8_u1_6734_wire(0) /=  '0') else IMC18_6554;
    -- logger for split-operator MUX_6745_inst flow-through 
    process(IMD10_6746) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6745_inst:flowthrough inputs: " & " BITSEL_u8_u1_6742_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6742_wire) & " IMC21_6578 = "& Convert_SLV_To_Hex_String(IMC21_6578) & " IMC20_6570 = "& Convert_SLV_To_Hex_String(IMC20_6570) & " outputs:" & " IMD10_6746= "  & Convert_SLV_To_Hex_String(IMD10_6746));
      --
    end process; 
    -- flow-through select operator MUX_6745_inst
    IMD10_6746 <= IMC21_6578 when (BITSEL_u8_u1_6742_wire(0) /=  '0') else IMC20_6570;
    -- logger for split-operator MUX_6753_inst flow-through 
    process(IMD11_6754) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6753_inst:flowthrough inputs: " & " BITSEL_u8_u1_6750_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6750_wire) & " IMC23_6594 = "& Convert_SLV_To_Hex_String(IMC23_6594) & " IMC22_6586 = "& Convert_SLV_To_Hex_String(IMC22_6586) & " outputs:" & " IMD11_6754= "  & Convert_SLV_To_Hex_String(IMD11_6754));
      --
    end process; 
    -- flow-through select operator MUX_6753_inst
    IMD11_6754 <= IMC23_6594 when (BITSEL_u8_u1_6750_wire(0) /=  '0') else IMC22_6586;
    -- logger for split-operator MUX_6761_inst flow-through 
    process(IMD12_6762) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6761_inst:flowthrough inputs: " & " BITSEL_u8_u1_6758_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6758_wire) & " IMC25_6610 = "& Convert_SLV_To_Hex_String(IMC25_6610) & " IMC24_6602 = "& Convert_SLV_To_Hex_String(IMC24_6602) & " outputs:" & " IMD12_6762= "  & Convert_SLV_To_Hex_String(IMD12_6762));
      --
    end process; 
    -- flow-through select operator MUX_6761_inst
    IMD12_6762 <= IMC25_6610 when (BITSEL_u8_u1_6758_wire(0) /=  '0') else IMC24_6602;
    -- logger for split-operator MUX_6769_inst flow-through 
    process(IMD13_6770) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6769_inst:flowthrough inputs: " & " BITSEL_u8_u1_6766_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6766_wire) & " IMC27_6626 = "& Convert_SLV_To_Hex_String(IMC27_6626) & " IMC26_6618 = "& Convert_SLV_To_Hex_String(IMC26_6618) & " outputs:" & " IMD13_6770= "  & Convert_SLV_To_Hex_String(IMD13_6770));
      --
    end process; 
    -- flow-through select operator MUX_6769_inst
    IMD13_6770 <= IMC27_6626 when (BITSEL_u8_u1_6766_wire(0) /=  '0') else IMC26_6618;
    -- logger for split-operator MUX_6777_inst flow-through 
    process(IMD14_6778) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6777_inst:flowthrough inputs: " & " BITSEL_u8_u1_6774_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6774_wire) & " IMC29_6642 = "& Convert_SLV_To_Hex_String(IMC29_6642) & " IMC28_6634 = "& Convert_SLV_To_Hex_String(IMC28_6634) & " outputs:" & " IMD14_6778= "  & Convert_SLV_To_Hex_String(IMD14_6778));
      --
    end process; 
    -- flow-through select operator MUX_6777_inst
    IMD14_6778 <= IMC29_6642 when (BITSEL_u8_u1_6774_wire(0) /=  '0') else IMC28_6634;
    -- logger for split-operator MUX_6785_inst flow-through 
    process(IMD15_6786) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6785_inst:flowthrough inputs: " & " BITSEL_u8_u1_6782_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6782_wire) & " IMC31_6658 = "& Convert_SLV_To_Hex_String(IMC31_6658) & " IMC30_6650 = "& Convert_SLV_To_Hex_String(IMC30_6650) & " outputs:" & " IMD15_6786= "  & Convert_SLV_To_Hex_String(IMD15_6786));
      --
    end process; 
    -- flow-through select operator MUX_6785_inst
    IMD15_6786 <= IMC31_6658 when (BITSEL_u8_u1_6782_wire(0) /=  '0') else IMC30_6650;
    -- logger for split-operator MUX_6793_inst flow-through 
    process(IME0_6794) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6793_inst:flowthrough inputs: " & " BITSEL_u8_u1_6790_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6790_wire) & " IMD1_6674 = "& Convert_SLV_To_Hex_String(IMD1_6674) & " IMD0_6666 = "& Convert_SLV_To_Hex_String(IMD0_6666) & " outputs:" & " IME0_6794= "  & Convert_SLV_To_Hex_String(IME0_6794));
      --
    end process; 
    -- flow-through select operator MUX_6793_inst
    IME0_6794 <= IMD1_6674 when (BITSEL_u8_u1_6790_wire(0) /=  '0') else IMD0_6666;
    -- logger for split-operator MUX_6801_inst flow-through 
    process(IME1_6802) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6801_inst:flowthrough inputs: " & " BITSEL_u8_u1_6798_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6798_wire) & " IMD3_6690 = "& Convert_SLV_To_Hex_String(IMD3_6690) & " IMD2_6682 = "& Convert_SLV_To_Hex_String(IMD2_6682) & " outputs:" & " IME1_6802= "  & Convert_SLV_To_Hex_String(IME1_6802));
      --
    end process; 
    -- flow-through select operator MUX_6801_inst
    IME1_6802 <= IMD3_6690 when (BITSEL_u8_u1_6798_wire(0) /=  '0') else IMD2_6682;
    -- logger for split-operator MUX_6809_inst flow-through 
    process(IME2_6810) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6809_inst:flowthrough inputs: " & " BITSEL_u8_u1_6806_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6806_wire) & " IMD5_6706 = "& Convert_SLV_To_Hex_String(IMD5_6706) & " IMD4_6698 = "& Convert_SLV_To_Hex_String(IMD4_6698) & " outputs:" & " IME2_6810= "  & Convert_SLV_To_Hex_String(IME2_6810));
      --
    end process; 
    -- flow-through select operator MUX_6809_inst
    IME2_6810 <= IMD5_6706 when (BITSEL_u8_u1_6806_wire(0) /=  '0') else IMD4_6698;
    -- logger for split-operator MUX_6817_inst flow-through 
    process(IME3_6818) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6817_inst:flowthrough inputs: " & " BITSEL_u8_u1_6814_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6814_wire) & " IMD7_6722 = "& Convert_SLV_To_Hex_String(IMD7_6722) & " IMD6_6714 = "& Convert_SLV_To_Hex_String(IMD6_6714) & " outputs:" & " IME3_6818= "  & Convert_SLV_To_Hex_String(IME3_6818));
      --
    end process; 
    -- flow-through select operator MUX_6817_inst
    IME3_6818 <= IMD7_6722 when (BITSEL_u8_u1_6814_wire(0) /=  '0') else IMD6_6714;
    -- logger for split-operator MUX_6825_inst flow-through 
    process(IME4_6826) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6825_inst:flowthrough inputs: " & " BITSEL_u8_u1_6822_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6822_wire) & " IMD9_6738 = "& Convert_SLV_To_Hex_String(IMD9_6738) & " IMD8_6730 = "& Convert_SLV_To_Hex_String(IMD8_6730) & " outputs:" & " IME4_6826= "  & Convert_SLV_To_Hex_String(IME4_6826));
      --
    end process; 
    -- flow-through select operator MUX_6825_inst
    IME4_6826 <= IMD9_6738 when (BITSEL_u8_u1_6822_wire(0) /=  '0') else IMD8_6730;
    -- logger for split-operator MUX_6833_inst flow-through 
    process(IME5_6834) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6833_inst:flowthrough inputs: " & " BITSEL_u8_u1_6830_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6830_wire) & " IMD11_6754 = "& Convert_SLV_To_Hex_String(IMD11_6754) & " IMD10_6746 = "& Convert_SLV_To_Hex_String(IMD10_6746) & " outputs:" & " IME5_6834= "  & Convert_SLV_To_Hex_String(IME5_6834));
      --
    end process; 
    -- flow-through select operator MUX_6833_inst
    IME5_6834 <= IMD11_6754 when (BITSEL_u8_u1_6830_wire(0) /=  '0') else IMD10_6746;
    -- logger for split-operator MUX_6841_inst flow-through 
    process(IME6_6842) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6841_inst:flowthrough inputs: " & " BITSEL_u8_u1_6838_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6838_wire) & " IMD13_6770 = "& Convert_SLV_To_Hex_String(IMD13_6770) & " IMD12_6762 = "& Convert_SLV_To_Hex_String(IMD12_6762) & " outputs:" & " IME6_6842= "  & Convert_SLV_To_Hex_String(IME6_6842));
      --
    end process; 
    -- flow-through select operator MUX_6841_inst
    IME6_6842 <= IMD13_6770 when (BITSEL_u8_u1_6838_wire(0) /=  '0') else IMD12_6762;
    -- logger for split-operator MUX_6849_inst flow-through 
    process(IME7_6850) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6849_inst:flowthrough inputs: " & " BITSEL_u8_u1_6846_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6846_wire) & " IMD15_6786 = "& Convert_SLV_To_Hex_String(IMD15_6786) & " IMD14_6778 = "& Convert_SLV_To_Hex_String(IMD14_6778) & " outputs:" & " IME7_6850= "  & Convert_SLV_To_Hex_String(IME7_6850));
      --
    end process; 
    -- flow-through select operator MUX_6849_inst
    IME7_6850 <= IMD15_6786 when (BITSEL_u8_u1_6846_wire(0) /=  '0') else IMD14_6778;
    -- logger for split-operator MUX_6857_inst flow-through 
    process(IMF0_6858) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6857_inst:flowthrough inputs: " & " BITSEL_u8_u1_6854_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6854_wire) & " IME1_6802 = "& Convert_SLV_To_Hex_String(IME1_6802) & " IME0_6794 = "& Convert_SLV_To_Hex_String(IME0_6794) & " outputs:" & " IMF0_6858= "  & Convert_SLV_To_Hex_String(IMF0_6858));
      --
    end process; 
    -- flow-through select operator MUX_6857_inst
    IMF0_6858 <= IME1_6802 when (BITSEL_u8_u1_6854_wire(0) /=  '0') else IME0_6794;
    -- logger for split-operator MUX_6865_inst flow-through 
    process(IMF1_6866) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6865_inst:flowthrough inputs: " & " BITSEL_u8_u1_6862_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6862_wire) & " IME3_6818 = "& Convert_SLV_To_Hex_String(IME3_6818) & " IME2_6810 = "& Convert_SLV_To_Hex_String(IME2_6810) & " outputs:" & " IMF1_6866= "  & Convert_SLV_To_Hex_String(IMF1_6866));
      --
    end process; 
    -- flow-through select operator MUX_6865_inst
    IMF1_6866 <= IME3_6818 when (BITSEL_u8_u1_6862_wire(0) /=  '0') else IME2_6810;
    -- logger for split-operator MUX_6873_inst flow-through 
    process(IMF2_6874) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6873_inst:flowthrough inputs: " & " BITSEL_u8_u1_6870_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6870_wire) & " IME5_6834 = "& Convert_SLV_To_Hex_String(IME5_6834) & " IME4_6826 = "& Convert_SLV_To_Hex_String(IME4_6826) & " outputs:" & " IMF2_6874= "  & Convert_SLV_To_Hex_String(IMF2_6874));
      --
    end process; 
    -- flow-through select operator MUX_6873_inst
    IMF2_6874 <= IME5_6834 when (BITSEL_u8_u1_6870_wire(0) /=  '0') else IME4_6826;
    -- logger for split-operator MUX_6881_inst flow-through 
    process(IMF3_6882) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6881_inst:flowthrough inputs: " & " BITSEL_u8_u1_6878_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6878_wire) & " IME7_6850 = "& Convert_SLV_To_Hex_String(IME7_6850) & " IME6_6842 = "& Convert_SLV_To_Hex_String(IME6_6842) & " outputs:" & " IMF3_6882= "  & Convert_SLV_To_Hex_String(IMF3_6882));
      --
    end process; 
    -- flow-through select operator MUX_6881_inst
    IMF3_6882 <= IME7_6850 when (BITSEL_u8_u1_6878_wire(0) /=  '0') else IME6_6842;
    -- logger for split-operator MUX_6889_inst flow-through 
    process(IMG0_6890) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6889_inst:flowthrough inputs: " & " BITSEL_u8_u1_6886_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6886_wire) & " IMF1_6866 = "& Convert_SLV_To_Hex_String(IMF1_6866) & " IMF0_6858 = "& Convert_SLV_To_Hex_String(IMF0_6858) & " outputs:" & " IMG0_6890= "  & Convert_SLV_To_Hex_String(IMG0_6890));
      --
    end process; 
    -- flow-through select operator MUX_6889_inst
    IMG0_6890 <= IMF1_6866 when (BITSEL_u8_u1_6886_wire(0) /=  '0') else IMF0_6858;
    -- logger for split-operator MUX_6897_inst flow-through 
    process(IMG1_6898) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6897_inst:flowthrough inputs: " & " BITSEL_u8_u1_6894_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6894_wire) & " IMF3_6882 = "& Convert_SLV_To_Hex_String(IMF3_6882) & " IMF2_6874 = "& Convert_SLV_To_Hex_String(IMF2_6874) & " outputs:" & " IMG1_6898= "  & Convert_SLV_To_Hex_String(IMG1_6898));
      --
    end process; 
    -- flow-through select operator MUX_6897_inst
    IMG1_6898 <= IMF3_6882 when (BITSEL_u8_u1_6894_wire(0) /=  '0') else IMF2_6874;
    -- logger for split-operator MUX_6905_inst flow-through 
    process(s_out_buffer) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:MUX_6905_inst:flowthrough inputs: " & " BITSEL_u8_u1_6902_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6902_wire) & " IMG1_6898 = "& Convert_SLV_To_Hex_String(IMG1_6898) & " IMG0_6890 = "& Convert_SLV_To_Hex_String(IMG0_6890) & " outputs:" & " s_out_buffer= "  & Convert_SLV_To_Hex_String(s_out_buffer));
      --
    end process; 
    -- flow-through select operator MUX_6905_inst
    s_out_buffer <= IMG1_6898 when (BITSEL_u8_u1_6902_wire(0) /=  '0') else IMG0_6890;
    -- logger for split-operator BITSEL_u8_u1_4614_inst flow-through 
    process(BITSEL_u8_u1_4614_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_4614_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4613_wire_constant = "& Convert_SLV_To_Hex_String(konst_4613_wire_constant) & " outputs:" & " BITSEL_u8_u1_4614_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4614_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4614_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4613_wire_constant, tmp_var);
      BITSEL_u8_u1_4614_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4624_inst flow-through 
    process(BITSEL_u8_u1_4624_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_4624_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4623_wire_constant = "& Convert_SLV_To_Hex_String(konst_4623_wire_constant) & " outputs:" & " BITSEL_u8_u1_4624_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4624_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4624_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4623_wire_constant, tmp_var);
      BITSEL_u8_u1_4624_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4634_inst flow-through 
    process(BITSEL_u8_u1_4634_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_4634_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4633_wire_constant = "& Convert_SLV_To_Hex_String(konst_4633_wire_constant) & " outputs:" & " BITSEL_u8_u1_4634_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4634_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4634_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4633_wire_constant, tmp_var);
      BITSEL_u8_u1_4634_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4644_inst flow-through 
    process(BITSEL_u8_u1_4644_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_4644_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4643_wire_constant = "& Convert_SLV_To_Hex_String(konst_4643_wire_constant) & " outputs:" & " BITSEL_u8_u1_4644_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4644_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4644_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4643_wire_constant, tmp_var);
      BITSEL_u8_u1_4644_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4654_inst flow-through 
    process(BITSEL_u8_u1_4654_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_4654_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4653_wire_constant = "& Convert_SLV_To_Hex_String(konst_4653_wire_constant) & " outputs:" & " BITSEL_u8_u1_4654_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4654_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4654_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4653_wire_constant, tmp_var);
      BITSEL_u8_u1_4654_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4664_inst flow-through 
    process(BITSEL_u8_u1_4664_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_4664_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4663_wire_constant = "& Convert_SLV_To_Hex_String(konst_4663_wire_constant) & " outputs:" & " BITSEL_u8_u1_4664_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4664_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4664_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4663_wire_constant, tmp_var);
      BITSEL_u8_u1_4664_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4674_inst flow-through 
    process(BITSEL_u8_u1_4674_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_4674_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4673_wire_constant = "& Convert_SLV_To_Hex_String(konst_4673_wire_constant) & " outputs:" & " BITSEL_u8_u1_4674_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4674_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4674_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4673_wire_constant, tmp_var);
      BITSEL_u8_u1_4674_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4684_inst flow-through 
    process(BITSEL_u8_u1_4684_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_4684_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4683_wire_constant = "& Convert_SLV_To_Hex_String(konst_4683_wire_constant) & " outputs:" & " BITSEL_u8_u1_4684_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4684_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4684_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4683_wire_constant, tmp_var);
      BITSEL_u8_u1_4684_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4694_inst flow-through 
    process(BITSEL_u8_u1_4694_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_4694_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4693_wire_constant = "& Convert_SLV_To_Hex_String(konst_4693_wire_constant) & " outputs:" & " BITSEL_u8_u1_4694_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4694_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4694_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4693_wire_constant, tmp_var);
      BITSEL_u8_u1_4694_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4704_inst flow-through 
    process(BITSEL_u8_u1_4704_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_4704_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4703_wire_constant = "& Convert_SLV_To_Hex_String(konst_4703_wire_constant) & " outputs:" & " BITSEL_u8_u1_4704_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4704_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4704_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4703_wire_constant, tmp_var);
      BITSEL_u8_u1_4704_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4714_inst flow-through 
    process(BITSEL_u8_u1_4714_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_4714_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4713_wire_constant = "& Convert_SLV_To_Hex_String(konst_4713_wire_constant) & " outputs:" & " BITSEL_u8_u1_4714_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4714_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4714_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4713_wire_constant, tmp_var);
      BITSEL_u8_u1_4714_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4724_inst flow-through 
    process(BITSEL_u8_u1_4724_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_4724_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4723_wire_constant = "& Convert_SLV_To_Hex_String(konst_4723_wire_constant) & " outputs:" & " BITSEL_u8_u1_4724_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4724_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4724_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4723_wire_constant, tmp_var);
      BITSEL_u8_u1_4724_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4734_inst flow-through 
    process(BITSEL_u8_u1_4734_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_4734_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4733_wire_constant = "& Convert_SLV_To_Hex_String(konst_4733_wire_constant) & " outputs:" & " BITSEL_u8_u1_4734_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4734_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4734_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4733_wire_constant, tmp_var);
      BITSEL_u8_u1_4734_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4744_inst flow-through 
    process(BITSEL_u8_u1_4744_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_4744_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4743_wire_constant = "& Convert_SLV_To_Hex_String(konst_4743_wire_constant) & " outputs:" & " BITSEL_u8_u1_4744_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4744_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4744_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4743_wire_constant, tmp_var);
      BITSEL_u8_u1_4744_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4754_inst flow-through 
    process(BITSEL_u8_u1_4754_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_4754_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4753_wire_constant = "& Convert_SLV_To_Hex_String(konst_4753_wire_constant) & " outputs:" & " BITSEL_u8_u1_4754_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4754_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4754_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4753_wire_constant, tmp_var);
      BITSEL_u8_u1_4754_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4764_inst flow-through 
    process(BITSEL_u8_u1_4764_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_4764_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4763_wire_constant = "& Convert_SLV_To_Hex_String(konst_4763_wire_constant) & " outputs:" & " BITSEL_u8_u1_4764_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4764_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4764_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4763_wire_constant, tmp_var);
      BITSEL_u8_u1_4764_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4774_inst flow-through 
    process(BITSEL_u8_u1_4774_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_4774_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4773_wire_constant = "& Convert_SLV_To_Hex_String(konst_4773_wire_constant) & " outputs:" & " BITSEL_u8_u1_4774_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4774_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4774_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4773_wire_constant, tmp_var);
      BITSEL_u8_u1_4774_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4784_inst flow-through 
    process(BITSEL_u8_u1_4784_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_4784_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4783_wire_constant = "& Convert_SLV_To_Hex_String(konst_4783_wire_constant) & " outputs:" & " BITSEL_u8_u1_4784_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4784_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4784_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4783_wire_constant, tmp_var);
      BITSEL_u8_u1_4784_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4794_inst flow-through 
    process(BITSEL_u8_u1_4794_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_4794_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4793_wire_constant = "& Convert_SLV_To_Hex_String(konst_4793_wire_constant) & " outputs:" & " BITSEL_u8_u1_4794_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4794_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4794_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4793_wire_constant, tmp_var);
      BITSEL_u8_u1_4794_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4804_inst flow-through 
    process(BITSEL_u8_u1_4804_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_4804_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4803_wire_constant = "& Convert_SLV_To_Hex_String(konst_4803_wire_constant) & " outputs:" & " BITSEL_u8_u1_4804_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4804_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4804_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4803_wire_constant, tmp_var);
      BITSEL_u8_u1_4804_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4814_inst flow-through 
    process(BITSEL_u8_u1_4814_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_4814_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4813_wire_constant = "& Convert_SLV_To_Hex_String(konst_4813_wire_constant) & " outputs:" & " BITSEL_u8_u1_4814_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4814_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4814_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4813_wire_constant, tmp_var);
      BITSEL_u8_u1_4814_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4824_inst flow-through 
    process(BITSEL_u8_u1_4824_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_4824_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4823_wire_constant = "& Convert_SLV_To_Hex_String(konst_4823_wire_constant) & " outputs:" & " BITSEL_u8_u1_4824_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4824_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4824_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4823_wire_constant, tmp_var);
      BITSEL_u8_u1_4824_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4834_inst flow-through 
    process(BITSEL_u8_u1_4834_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_4834_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4833_wire_constant = "& Convert_SLV_To_Hex_String(konst_4833_wire_constant) & " outputs:" & " BITSEL_u8_u1_4834_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4834_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4834_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4833_wire_constant, tmp_var);
      BITSEL_u8_u1_4834_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4844_inst flow-through 
    process(BITSEL_u8_u1_4844_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_4844_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4843_wire_constant = "& Convert_SLV_To_Hex_String(konst_4843_wire_constant) & " outputs:" & " BITSEL_u8_u1_4844_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4844_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4844_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4843_wire_constant, tmp_var);
      BITSEL_u8_u1_4844_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4854_inst flow-through 
    process(BITSEL_u8_u1_4854_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_4854_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4853_wire_constant = "& Convert_SLV_To_Hex_String(konst_4853_wire_constant) & " outputs:" & " BITSEL_u8_u1_4854_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4854_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4854_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4853_wire_constant, tmp_var);
      BITSEL_u8_u1_4854_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4864_inst flow-through 
    process(BITSEL_u8_u1_4864_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_4864_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4863_wire_constant = "& Convert_SLV_To_Hex_String(konst_4863_wire_constant) & " outputs:" & " BITSEL_u8_u1_4864_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4864_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4864_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4863_wire_constant, tmp_var);
      BITSEL_u8_u1_4864_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4874_inst flow-through 
    process(BITSEL_u8_u1_4874_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_4874_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4873_wire_constant = "& Convert_SLV_To_Hex_String(konst_4873_wire_constant) & " outputs:" & " BITSEL_u8_u1_4874_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4874_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4874_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4873_wire_constant, tmp_var);
      BITSEL_u8_u1_4874_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4884_inst flow-through 
    process(BITSEL_u8_u1_4884_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_4884_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4883_wire_constant = "& Convert_SLV_To_Hex_String(konst_4883_wire_constant) & " outputs:" & " BITSEL_u8_u1_4884_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4884_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4884_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4883_wire_constant, tmp_var);
      BITSEL_u8_u1_4884_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4894_inst flow-through 
    process(BITSEL_u8_u1_4894_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_4894_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4893_wire_constant = "& Convert_SLV_To_Hex_String(konst_4893_wire_constant) & " outputs:" & " BITSEL_u8_u1_4894_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4894_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4894_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4893_wire_constant, tmp_var);
      BITSEL_u8_u1_4894_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4904_inst flow-through 
    process(BITSEL_u8_u1_4904_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_4904_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4903_wire_constant = "& Convert_SLV_To_Hex_String(konst_4903_wire_constant) & " outputs:" & " BITSEL_u8_u1_4904_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4904_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4904_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4903_wire_constant, tmp_var);
      BITSEL_u8_u1_4904_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4914_inst flow-through 
    process(BITSEL_u8_u1_4914_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_4914_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4913_wire_constant = "& Convert_SLV_To_Hex_String(konst_4913_wire_constant) & " outputs:" & " BITSEL_u8_u1_4914_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4914_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4914_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4913_wire_constant, tmp_var);
      BITSEL_u8_u1_4914_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4924_inst flow-through 
    process(BITSEL_u8_u1_4924_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_4924_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4923_wire_constant = "& Convert_SLV_To_Hex_String(konst_4923_wire_constant) & " outputs:" & " BITSEL_u8_u1_4924_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4924_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4924_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4923_wire_constant, tmp_var);
      BITSEL_u8_u1_4924_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4934_inst flow-through 
    process(BITSEL_u8_u1_4934_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_4934_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4933_wire_constant = "& Convert_SLV_To_Hex_String(konst_4933_wire_constant) & " outputs:" & " BITSEL_u8_u1_4934_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4934_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4934_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4933_wire_constant, tmp_var);
      BITSEL_u8_u1_4934_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4944_inst flow-through 
    process(BITSEL_u8_u1_4944_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_4944_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4943_wire_constant = "& Convert_SLV_To_Hex_String(konst_4943_wire_constant) & " outputs:" & " BITSEL_u8_u1_4944_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4944_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4944_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4943_wire_constant, tmp_var);
      BITSEL_u8_u1_4944_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4954_inst flow-through 
    process(BITSEL_u8_u1_4954_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_4954_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4953_wire_constant = "& Convert_SLV_To_Hex_String(konst_4953_wire_constant) & " outputs:" & " BITSEL_u8_u1_4954_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4954_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4954_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4953_wire_constant, tmp_var);
      BITSEL_u8_u1_4954_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4964_inst flow-through 
    process(BITSEL_u8_u1_4964_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_4964_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4963_wire_constant = "& Convert_SLV_To_Hex_String(konst_4963_wire_constant) & " outputs:" & " BITSEL_u8_u1_4964_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4964_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4964_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4963_wire_constant, tmp_var);
      BITSEL_u8_u1_4964_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4974_inst flow-through 
    process(BITSEL_u8_u1_4974_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_4974_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4973_wire_constant = "& Convert_SLV_To_Hex_String(konst_4973_wire_constant) & " outputs:" & " BITSEL_u8_u1_4974_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4974_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4974_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4973_wire_constant, tmp_var);
      BITSEL_u8_u1_4974_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4984_inst flow-through 
    process(BITSEL_u8_u1_4984_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_4984_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4983_wire_constant = "& Convert_SLV_To_Hex_String(konst_4983_wire_constant) & " outputs:" & " BITSEL_u8_u1_4984_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4984_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4984_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4983_wire_constant, tmp_var);
      BITSEL_u8_u1_4984_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_4994_inst flow-through 
    process(BITSEL_u8_u1_4994_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_4994_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_4993_wire_constant = "& Convert_SLV_To_Hex_String(konst_4993_wire_constant) & " outputs:" & " BITSEL_u8_u1_4994_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_4994_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_4994_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4993_wire_constant, tmp_var);
      BITSEL_u8_u1_4994_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_5004_inst flow-through 
    process(BITSEL_u8_u1_5004_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_5004_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_5003_wire_constant = "& Convert_SLV_To_Hex_String(konst_5003_wire_constant) & " outputs:" & " BITSEL_u8_u1_5004_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_5004_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_5004_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5003_wire_constant, tmp_var);
      BITSEL_u8_u1_5004_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_5014_inst flow-through 
    process(BITSEL_u8_u1_5014_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_5014_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_5013_wire_constant = "& Convert_SLV_To_Hex_String(konst_5013_wire_constant) & " outputs:" & " BITSEL_u8_u1_5014_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_5014_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_5014_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5013_wire_constant, tmp_var);
      BITSEL_u8_u1_5014_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_5024_inst flow-through 
    process(BITSEL_u8_u1_5024_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_5024_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_5023_wire_constant = "& Convert_SLV_To_Hex_String(konst_5023_wire_constant) & " outputs:" & " BITSEL_u8_u1_5024_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_5024_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_5024_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5023_wire_constant, tmp_var);
      BITSEL_u8_u1_5024_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_5034_inst flow-through 
    process(BITSEL_u8_u1_5034_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_5034_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_5033_wire_constant = "& Convert_SLV_To_Hex_String(konst_5033_wire_constant) & " outputs:" & " BITSEL_u8_u1_5034_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_5034_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_5034_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5033_wire_constant, tmp_var);
      BITSEL_u8_u1_5034_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_5044_inst flow-through 
    process(BITSEL_u8_u1_5044_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_5044_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_5043_wire_constant = "& Convert_SLV_To_Hex_String(konst_5043_wire_constant) & " outputs:" & " BITSEL_u8_u1_5044_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_5044_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_5044_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5043_wire_constant, tmp_var);
      BITSEL_u8_u1_5044_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_5054_inst flow-through 
    process(BITSEL_u8_u1_5054_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_5054_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_5053_wire_constant = "& Convert_SLV_To_Hex_String(konst_5053_wire_constant) & " outputs:" & " BITSEL_u8_u1_5054_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_5054_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_5054_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5053_wire_constant, tmp_var);
      BITSEL_u8_u1_5054_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_5064_inst flow-through 
    process(BITSEL_u8_u1_5064_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_5064_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_5063_wire_constant = "& Convert_SLV_To_Hex_String(konst_5063_wire_constant) & " outputs:" & " BITSEL_u8_u1_5064_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_5064_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_5064_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5063_wire_constant, tmp_var);
      BITSEL_u8_u1_5064_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_5074_inst flow-through 
    process(BITSEL_u8_u1_5074_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_5074_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_5073_wire_constant = "& Convert_SLV_To_Hex_String(konst_5073_wire_constant) & " outputs:" & " BITSEL_u8_u1_5074_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_5074_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_5074_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5073_wire_constant, tmp_var);
      BITSEL_u8_u1_5074_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_5084_inst flow-through 
    process(BITSEL_u8_u1_5084_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_5084_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_5083_wire_constant = "& Convert_SLV_To_Hex_String(konst_5083_wire_constant) & " outputs:" & " BITSEL_u8_u1_5084_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_5084_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_5084_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5083_wire_constant, tmp_var);
      BITSEL_u8_u1_5084_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_5094_inst flow-through 
    process(BITSEL_u8_u1_5094_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_5094_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_5093_wire_constant = "& Convert_SLV_To_Hex_String(konst_5093_wire_constant) & " outputs:" & " BITSEL_u8_u1_5094_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_5094_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_5094_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5093_wire_constant, tmp_var);
      BITSEL_u8_u1_5094_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_5104_inst flow-through 
    process(BITSEL_u8_u1_5104_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_5104_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_5103_wire_constant = "& Convert_SLV_To_Hex_String(konst_5103_wire_constant) & " outputs:" & " BITSEL_u8_u1_5104_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_5104_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_5104_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5103_wire_constant, tmp_var);
      BITSEL_u8_u1_5104_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_5114_inst flow-through 
    process(BITSEL_u8_u1_5114_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_5114_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_5113_wire_constant = "& Convert_SLV_To_Hex_String(konst_5113_wire_constant) & " outputs:" & " BITSEL_u8_u1_5114_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_5114_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_5114_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5113_wire_constant, tmp_var);
      BITSEL_u8_u1_5114_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_5124_inst flow-through 
    process(BITSEL_u8_u1_5124_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_5124_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_5123_wire_constant = "& Convert_SLV_To_Hex_String(konst_5123_wire_constant) & " outputs:" & " BITSEL_u8_u1_5124_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_5124_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_5124_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5123_wire_constant, tmp_var);
      BITSEL_u8_u1_5124_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_5134_inst flow-through 
    process(BITSEL_u8_u1_5134_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_5134_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_5133_wire_constant = "& Convert_SLV_To_Hex_String(konst_5133_wire_constant) & " outputs:" & " BITSEL_u8_u1_5134_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_5134_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_5134_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5133_wire_constant, tmp_var);
      BITSEL_u8_u1_5134_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_5144_inst flow-through 
    process(BITSEL_u8_u1_5144_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_5144_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_5143_wire_constant = "& Convert_SLV_To_Hex_String(konst_5143_wire_constant) & " outputs:" & " BITSEL_u8_u1_5144_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_5144_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_5144_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5143_wire_constant, tmp_var);
      BITSEL_u8_u1_5144_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_5154_inst flow-through 
    process(BITSEL_u8_u1_5154_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_5154_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_5153_wire_constant = "& Convert_SLV_To_Hex_String(konst_5153_wire_constant) & " outputs:" & " BITSEL_u8_u1_5154_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_5154_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_5154_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5153_wire_constant, tmp_var);
      BITSEL_u8_u1_5154_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_5164_inst flow-through 
    process(BITSEL_u8_u1_5164_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_5164_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_5163_wire_constant = "& Convert_SLV_To_Hex_String(konst_5163_wire_constant) & " outputs:" & " BITSEL_u8_u1_5164_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_5164_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_5164_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5163_wire_constant, tmp_var);
      BITSEL_u8_u1_5164_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_5174_inst flow-through 
    process(BITSEL_u8_u1_5174_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_5174_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_5173_wire_constant = "& Convert_SLV_To_Hex_String(konst_5173_wire_constant) & " outputs:" & " BITSEL_u8_u1_5174_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_5174_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_5174_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5173_wire_constant, tmp_var);
      BITSEL_u8_u1_5174_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_5184_inst flow-through 
    process(BITSEL_u8_u1_5184_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_5184_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_5183_wire_constant = "& Convert_SLV_To_Hex_String(konst_5183_wire_constant) & " outputs:" & " BITSEL_u8_u1_5184_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_5184_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_5184_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5183_wire_constant, tmp_var);
      BITSEL_u8_u1_5184_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_5194_inst flow-through 
    process(BITSEL_u8_u1_5194_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_5194_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_5193_wire_constant = "& Convert_SLV_To_Hex_String(konst_5193_wire_constant) & " outputs:" & " BITSEL_u8_u1_5194_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_5194_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_5194_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5193_wire_constant, tmp_var);
      BITSEL_u8_u1_5194_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_5204_inst flow-through 
    process(BITSEL_u8_u1_5204_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_5204_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_5203_wire_constant = "& Convert_SLV_To_Hex_String(konst_5203_wire_constant) & " outputs:" & " BITSEL_u8_u1_5204_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_5204_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_5204_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5203_wire_constant, tmp_var);
      BITSEL_u8_u1_5204_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_5214_inst flow-through 
    process(BITSEL_u8_u1_5214_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_5214_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_5213_wire_constant = "& Convert_SLV_To_Hex_String(konst_5213_wire_constant) & " outputs:" & " BITSEL_u8_u1_5214_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_5214_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_5214_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5213_wire_constant, tmp_var);
      BITSEL_u8_u1_5214_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_5224_inst flow-through 
    process(BITSEL_u8_u1_5224_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_5224_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_5223_wire_constant = "& Convert_SLV_To_Hex_String(konst_5223_wire_constant) & " outputs:" & " BITSEL_u8_u1_5224_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_5224_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_5224_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5223_wire_constant, tmp_var);
      BITSEL_u8_u1_5224_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_5234_inst flow-through 
    process(BITSEL_u8_u1_5234_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_5234_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_5233_wire_constant = "& Convert_SLV_To_Hex_String(konst_5233_wire_constant) & " outputs:" & " BITSEL_u8_u1_5234_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_5234_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_5234_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5233_wire_constant, tmp_var);
      BITSEL_u8_u1_5234_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_5244_inst flow-through 
    process(BITSEL_u8_u1_5244_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_5244_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_5243_wire_constant = "& Convert_SLV_To_Hex_String(konst_5243_wire_constant) & " outputs:" & " BITSEL_u8_u1_5244_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_5244_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_5244_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5243_wire_constant, tmp_var);
      BITSEL_u8_u1_5244_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_5254_inst flow-through 
    process(BITSEL_u8_u1_5254_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_5254_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_5253_wire_constant = "& Convert_SLV_To_Hex_String(konst_5253_wire_constant) & " outputs:" & " BITSEL_u8_u1_5254_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_5254_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_5254_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5253_wire_constant, tmp_var);
      BITSEL_u8_u1_5254_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_5264_inst flow-through 
    process(BITSEL_u8_u1_5264_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_5264_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_5263_wire_constant = "& Convert_SLV_To_Hex_String(konst_5263_wire_constant) & " outputs:" & " BITSEL_u8_u1_5264_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_5264_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_5264_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5263_wire_constant, tmp_var);
      BITSEL_u8_u1_5264_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_5274_inst flow-through 
    process(BITSEL_u8_u1_5274_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_5274_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_5273_wire_constant = "& Convert_SLV_To_Hex_String(konst_5273_wire_constant) & " outputs:" & " BITSEL_u8_u1_5274_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_5274_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_5274_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5273_wire_constant, tmp_var);
      BITSEL_u8_u1_5274_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_5284_inst flow-through 
    process(BITSEL_u8_u1_5284_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_5284_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_5283_wire_constant = "& Convert_SLV_To_Hex_String(konst_5283_wire_constant) & " outputs:" & " BITSEL_u8_u1_5284_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_5284_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_5284_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5283_wire_constant, tmp_var);
      BITSEL_u8_u1_5284_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_5294_inst flow-through 
    process(BITSEL_u8_u1_5294_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_5294_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_5293_wire_constant = "& Convert_SLV_To_Hex_String(konst_5293_wire_constant) & " outputs:" & " BITSEL_u8_u1_5294_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_5294_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_5294_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5293_wire_constant, tmp_var);
      BITSEL_u8_u1_5294_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_5304_inst flow-through 
    process(BITSEL_u8_u1_5304_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_5304_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_5303_wire_constant = "& Convert_SLV_To_Hex_String(konst_5303_wire_constant) & " outputs:" & " BITSEL_u8_u1_5304_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_5304_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_5304_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5303_wire_constant, tmp_var);
      BITSEL_u8_u1_5304_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_5314_inst flow-through 
    process(BITSEL_u8_u1_5314_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_5314_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_5313_wire_constant = "& Convert_SLV_To_Hex_String(konst_5313_wire_constant) & " outputs:" & " BITSEL_u8_u1_5314_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_5314_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_5314_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5313_wire_constant, tmp_var);
      BITSEL_u8_u1_5314_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_5324_inst flow-through 
    process(BITSEL_u8_u1_5324_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_5324_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_5323_wire_constant = "& Convert_SLV_To_Hex_String(konst_5323_wire_constant) & " outputs:" & " BITSEL_u8_u1_5324_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_5324_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_5324_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5323_wire_constant, tmp_var);
      BITSEL_u8_u1_5324_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_5334_inst flow-through 
    process(BITSEL_u8_u1_5334_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_5334_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_5333_wire_constant = "& Convert_SLV_To_Hex_String(konst_5333_wire_constant) & " outputs:" & " BITSEL_u8_u1_5334_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_5334_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_5334_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5333_wire_constant, tmp_var);
      BITSEL_u8_u1_5334_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_5344_inst flow-through 
    process(BITSEL_u8_u1_5344_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_5344_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_5343_wire_constant = "& Convert_SLV_To_Hex_String(konst_5343_wire_constant) & " outputs:" & " BITSEL_u8_u1_5344_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_5344_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_5344_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5343_wire_constant, tmp_var);
      BITSEL_u8_u1_5344_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_5354_inst flow-through 
    process(BITSEL_u8_u1_5354_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_5354_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_5353_wire_constant = "& Convert_SLV_To_Hex_String(konst_5353_wire_constant) & " outputs:" & " BITSEL_u8_u1_5354_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_5354_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_5354_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5353_wire_constant, tmp_var);
      BITSEL_u8_u1_5354_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_5364_inst flow-through 
    process(BITSEL_u8_u1_5364_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_5364_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_5363_wire_constant = "& Convert_SLV_To_Hex_String(konst_5363_wire_constant) & " outputs:" & " BITSEL_u8_u1_5364_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_5364_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_5364_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5363_wire_constant, tmp_var);
      BITSEL_u8_u1_5364_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_5374_inst flow-through 
    process(BITSEL_u8_u1_5374_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_5374_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_5373_wire_constant = "& Convert_SLV_To_Hex_String(konst_5373_wire_constant) & " outputs:" & " BITSEL_u8_u1_5374_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_5374_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_5374_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5373_wire_constant, tmp_var);
      BITSEL_u8_u1_5374_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_5384_inst flow-through 
    process(BITSEL_u8_u1_5384_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_5384_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_5383_wire_constant = "& Convert_SLV_To_Hex_String(konst_5383_wire_constant) & " outputs:" & " BITSEL_u8_u1_5384_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_5384_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_5384_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5383_wire_constant, tmp_var);
      BITSEL_u8_u1_5384_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_5394_inst flow-through 
    process(BITSEL_u8_u1_5394_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_5394_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_5393_wire_constant = "& Convert_SLV_To_Hex_String(konst_5393_wire_constant) & " outputs:" & " BITSEL_u8_u1_5394_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_5394_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_5394_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5393_wire_constant, tmp_var);
      BITSEL_u8_u1_5394_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_5404_inst flow-through 
    process(BITSEL_u8_u1_5404_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_5404_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_5403_wire_constant = "& Convert_SLV_To_Hex_String(konst_5403_wire_constant) & " outputs:" & " BITSEL_u8_u1_5404_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_5404_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_5404_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5403_wire_constant, tmp_var);
      BITSEL_u8_u1_5404_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_5414_inst flow-through 
    process(BITSEL_u8_u1_5414_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_5414_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_5413_wire_constant = "& Convert_SLV_To_Hex_String(konst_5413_wire_constant) & " outputs:" & " BITSEL_u8_u1_5414_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_5414_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_5414_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5413_wire_constant, tmp_var);
      BITSEL_u8_u1_5414_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_5424_inst flow-through 
    process(BITSEL_u8_u1_5424_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_5424_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_5423_wire_constant = "& Convert_SLV_To_Hex_String(konst_5423_wire_constant) & " outputs:" & " BITSEL_u8_u1_5424_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_5424_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_5424_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5423_wire_constant, tmp_var);
      BITSEL_u8_u1_5424_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_5434_inst flow-through 
    process(BITSEL_u8_u1_5434_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_5434_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_5433_wire_constant = "& Convert_SLV_To_Hex_String(konst_5433_wire_constant) & " outputs:" & " BITSEL_u8_u1_5434_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_5434_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_5434_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5433_wire_constant, tmp_var);
      BITSEL_u8_u1_5434_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_5444_inst flow-through 
    process(BITSEL_u8_u1_5444_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_5444_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_5443_wire_constant = "& Convert_SLV_To_Hex_String(konst_5443_wire_constant) & " outputs:" & " BITSEL_u8_u1_5444_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_5444_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_5444_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5443_wire_constant, tmp_var);
      BITSEL_u8_u1_5444_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_5454_inst flow-through 
    process(BITSEL_u8_u1_5454_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_5454_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_5453_wire_constant = "& Convert_SLV_To_Hex_String(konst_5453_wire_constant) & " outputs:" & " BITSEL_u8_u1_5454_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_5454_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_5454_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5453_wire_constant, tmp_var);
      BITSEL_u8_u1_5454_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_5464_inst flow-through 
    process(BITSEL_u8_u1_5464_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_5464_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_5463_wire_constant = "& Convert_SLV_To_Hex_String(konst_5463_wire_constant) & " outputs:" & " BITSEL_u8_u1_5464_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_5464_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_5464_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5463_wire_constant, tmp_var);
      BITSEL_u8_u1_5464_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_5474_inst flow-through 
    process(BITSEL_u8_u1_5474_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_5474_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_5473_wire_constant = "& Convert_SLV_To_Hex_String(konst_5473_wire_constant) & " outputs:" & " BITSEL_u8_u1_5474_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_5474_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_5474_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5473_wire_constant, tmp_var);
      BITSEL_u8_u1_5474_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_5484_inst flow-through 
    process(BITSEL_u8_u1_5484_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_5484_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_5483_wire_constant = "& Convert_SLV_To_Hex_String(konst_5483_wire_constant) & " outputs:" & " BITSEL_u8_u1_5484_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_5484_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_5484_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5483_wire_constant, tmp_var);
      BITSEL_u8_u1_5484_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_5494_inst flow-through 
    process(BITSEL_u8_u1_5494_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_5494_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_5493_wire_constant = "& Convert_SLV_To_Hex_String(konst_5493_wire_constant) & " outputs:" & " BITSEL_u8_u1_5494_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_5494_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_5494_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5493_wire_constant, tmp_var);
      BITSEL_u8_u1_5494_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_5504_inst flow-through 
    process(BITSEL_u8_u1_5504_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_5504_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_5503_wire_constant = "& Convert_SLV_To_Hex_String(konst_5503_wire_constant) & " outputs:" & " BITSEL_u8_u1_5504_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_5504_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_5504_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5503_wire_constant, tmp_var);
      BITSEL_u8_u1_5504_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_5514_inst flow-through 
    process(BITSEL_u8_u1_5514_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_5514_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_5513_wire_constant = "& Convert_SLV_To_Hex_String(konst_5513_wire_constant) & " outputs:" & " BITSEL_u8_u1_5514_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_5514_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_5514_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5513_wire_constant, tmp_var);
      BITSEL_u8_u1_5514_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_5524_inst flow-through 
    process(BITSEL_u8_u1_5524_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_5524_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_5523_wire_constant = "& Convert_SLV_To_Hex_String(konst_5523_wire_constant) & " outputs:" & " BITSEL_u8_u1_5524_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_5524_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_5524_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5523_wire_constant, tmp_var);
      BITSEL_u8_u1_5524_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_5534_inst flow-through 
    process(BITSEL_u8_u1_5534_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_5534_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_5533_wire_constant = "& Convert_SLV_To_Hex_String(konst_5533_wire_constant) & " outputs:" & " BITSEL_u8_u1_5534_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_5534_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_5534_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5533_wire_constant, tmp_var);
      BITSEL_u8_u1_5534_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_5544_inst flow-through 
    process(BITSEL_u8_u1_5544_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_5544_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_5543_wire_constant = "& Convert_SLV_To_Hex_String(konst_5543_wire_constant) & " outputs:" & " BITSEL_u8_u1_5544_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_5544_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_5544_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5543_wire_constant, tmp_var);
      BITSEL_u8_u1_5544_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_5554_inst flow-through 
    process(BITSEL_u8_u1_5554_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_5554_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_5553_wire_constant = "& Convert_SLV_To_Hex_String(konst_5553_wire_constant) & " outputs:" & " BITSEL_u8_u1_5554_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_5554_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_5554_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5553_wire_constant, tmp_var);
      BITSEL_u8_u1_5554_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_5564_inst flow-through 
    process(BITSEL_u8_u1_5564_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_5564_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_5563_wire_constant = "& Convert_SLV_To_Hex_String(konst_5563_wire_constant) & " outputs:" & " BITSEL_u8_u1_5564_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_5564_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_5564_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5563_wire_constant, tmp_var);
      BITSEL_u8_u1_5564_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_5574_inst flow-through 
    process(BITSEL_u8_u1_5574_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_5574_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_5573_wire_constant = "& Convert_SLV_To_Hex_String(konst_5573_wire_constant) & " outputs:" & " BITSEL_u8_u1_5574_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_5574_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_5574_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5573_wire_constant, tmp_var);
      BITSEL_u8_u1_5574_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_5584_inst flow-through 
    process(BITSEL_u8_u1_5584_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_5584_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_5583_wire_constant = "& Convert_SLV_To_Hex_String(konst_5583_wire_constant) & " outputs:" & " BITSEL_u8_u1_5584_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_5584_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_5584_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5583_wire_constant, tmp_var);
      BITSEL_u8_u1_5584_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_5594_inst flow-through 
    process(BITSEL_u8_u1_5594_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_5594_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_5593_wire_constant = "& Convert_SLV_To_Hex_String(konst_5593_wire_constant) & " outputs:" & " BITSEL_u8_u1_5594_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_5594_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_5594_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5593_wire_constant, tmp_var);
      BITSEL_u8_u1_5594_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_5604_inst flow-through 
    process(BITSEL_u8_u1_5604_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_5604_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_5603_wire_constant = "& Convert_SLV_To_Hex_String(konst_5603_wire_constant) & " outputs:" & " BITSEL_u8_u1_5604_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_5604_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_5604_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5603_wire_constant, tmp_var);
      BITSEL_u8_u1_5604_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_5614_inst flow-through 
    process(BITSEL_u8_u1_5614_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_5614_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_5613_wire_constant = "& Convert_SLV_To_Hex_String(konst_5613_wire_constant) & " outputs:" & " BITSEL_u8_u1_5614_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_5614_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_5614_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5613_wire_constant, tmp_var);
      BITSEL_u8_u1_5614_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_5624_inst flow-through 
    process(BITSEL_u8_u1_5624_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_5624_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_5623_wire_constant = "& Convert_SLV_To_Hex_String(konst_5623_wire_constant) & " outputs:" & " BITSEL_u8_u1_5624_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_5624_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_5624_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5623_wire_constant, tmp_var);
      BITSEL_u8_u1_5624_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_5634_inst flow-through 
    process(BITSEL_u8_u1_5634_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_5634_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_5633_wire_constant = "& Convert_SLV_To_Hex_String(konst_5633_wire_constant) & " outputs:" & " BITSEL_u8_u1_5634_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_5634_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_5634_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5633_wire_constant, tmp_var);
      BITSEL_u8_u1_5634_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_5644_inst flow-through 
    process(BITSEL_u8_u1_5644_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_5644_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_5643_wire_constant = "& Convert_SLV_To_Hex_String(konst_5643_wire_constant) & " outputs:" & " BITSEL_u8_u1_5644_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_5644_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_5644_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5643_wire_constant, tmp_var);
      BITSEL_u8_u1_5644_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_5654_inst flow-through 
    process(BITSEL_u8_u1_5654_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_5654_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_5653_wire_constant = "& Convert_SLV_To_Hex_String(konst_5653_wire_constant) & " outputs:" & " BITSEL_u8_u1_5654_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_5654_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_5654_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5653_wire_constant, tmp_var);
      BITSEL_u8_u1_5654_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_5664_inst flow-through 
    process(BITSEL_u8_u1_5664_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_5664_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_5663_wire_constant = "& Convert_SLV_To_Hex_String(konst_5663_wire_constant) & " outputs:" & " BITSEL_u8_u1_5664_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_5664_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_5664_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5663_wire_constant, tmp_var);
      BITSEL_u8_u1_5664_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_5674_inst flow-through 
    process(BITSEL_u8_u1_5674_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_5674_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_5673_wire_constant = "& Convert_SLV_To_Hex_String(konst_5673_wire_constant) & " outputs:" & " BITSEL_u8_u1_5674_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_5674_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_5674_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5673_wire_constant, tmp_var);
      BITSEL_u8_u1_5674_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_5684_inst flow-through 
    process(BITSEL_u8_u1_5684_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_5684_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_5683_wire_constant = "& Convert_SLV_To_Hex_String(konst_5683_wire_constant) & " outputs:" & " BITSEL_u8_u1_5684_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_5684_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_5684_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5683_wire_constant, tmp_var);
      BITSEL_u8_u1_5684_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_5694_inst flow-through 
    process(BITSEL_u8_u1_5694_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_5694_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_5693_wire_constant = "& Convert_SLV_To_Hex_String(konst_5693_wire_constant) & " outputs:" & " BITSEL_u8_u1_5694_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_5694_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_5694_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5693_wire_constant, tmp_var);
      BITSEL_u8_u1_5694_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_5704_inst flow-through 
    process(BITSEL_u8_u1_5704_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_5704_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_5703_wire_constant = "& Convert_SLV_To_Hex_String(konst_5703_wire_constant) & " outputs:" & " BITSEL_u8_u1_5704_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_5704_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_5704_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5703_wire_constant, tmp_var);
      BITSEL_u8_u1_5704_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_5714_inst flow-through 
    process(BITSEL_u8_u1_5714_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_5714_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_5713_wire_constant = "& Convert_SLV_To_Hex_String(konst_5713_wire_constant) & " outputs:" & " BITSEL_u8_u1_5714_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_5714_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_5714_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5713_wire_constant, tmp_var);
      BITSEL_u8_u1_5714_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_5724_inst flow-through 
    process(BITSEL_u8_u1_5724_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_5724_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_5723_wire_constant = "& Convert_SLV_To_Hex_String(konst_5723_wire_constant) & " outputs:" & " BITSEL_u8_u1_5724_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_5724_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_5724_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5723_wire_constant, tmp_var);
      BITSEL_u8_u1_5724_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_5734_inst flow-through 
    process(BITSEL_u8_u1_5734_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_5734_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_5733_wire_constant = "& Convert_SLV_To_Hex_String(konst_5733_wire_constant) & " outputs:" & " BITSEL_u8_u1_5734_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_5734_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_5734_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5733_wire_constant, tmp_var);
      BITSEL_u8_u1_5734_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_5744_inst flow-through 
    process(BITSEL_u8_u1_5744_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_5744_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_5743_wire_constant = "& Convert_SLV_To_Hex_String(konst_5743_wire_constant) & " outputs:" & " BITSEL_u8_u1_5744_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_5744_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_5744_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5743_wire_constant, tmp_var);
      BITSEL_u8_u1_5744_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_5754_inst flow-through 
    process(BITSEL_u8_u1_5754_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_5754_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_5753_wire_constant = "& Convert_SLV_To_Hex_String(konst_5753_wire_constant) & " outputs:" & " BITSEL_u8_u1_5754_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_5754_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_5754_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5753_wire_constant, tmp_var);
      BITSEL_u8_u1_5754_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_5764_inst flow-through 
    process(BITSEL_u8_u1_5764_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_5764_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_5763_wire_constant = "& Convert_SLV_To_Hex_String(konst_5763_wire_constant) & " outputs:" & " BITSEL_u8_u1_5764_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_5764_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_5764_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5763_wire_constant, tmp_var);
      BITSEL_u8_u1_5764_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_5774_inst flow-through 
    process(BITSEL_u8_u1_5774_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_5774_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_5773_wire_constant = "& Convert_SLV_To_Hex_String(konst_5773_wire_constant) & " outputs:" & " BITSEL_u8_u1_5774_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_5774_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_5774_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5773_wire_constant, tmp_var);
      BITSEL_u8_u1_5774_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_5784_inst flow-through 
    process(BITSEL_u8_u1_5784_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_5784_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_5783_wire_constant = "& Convert_SLV_To_Hex_String(konst_5783_wire_constant) & " outputs:" & " BITSEL_u8_u1_5784_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_5784_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_5784_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5783_wire_constant, tmp_var);
      BITSEL_u8_u1_5784_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_5794_inst flow-through 
    process(BITSEL_u8_u1_5794_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_5794_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_5793_wire_constant = "& Convert_SLV_To_Hex_String(konst_5793_wire_constant) & " outputs:" & " BITSEL_u8_u1_5794_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_5794_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_5794_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5793_wire_constant, tmp_var);
      BITSEL_u8_u1_5794_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_5804_inst flow-through 
    process(BITSEL_u8_u1_5804_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_5804_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_5803_wire_constant = "& Convert_SLV_To_Hex_String(konst_5803_wire_constant) & " outputs:" & " BITSEL_u8_u1_5804_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_5804_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_5804_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5803_wire_constant, tmp_var);
      BITSEL_u8_u1_5804_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_5814_inst flow-through 
    process(BITSEL_u8_u1_5814_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_5814_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_5813_wire_constant = "& Convert_SLV_To_Hex_String(konst_5813_wire_constant) & " outputs:" & " BITSEL_u8_u1_5814_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_5814_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_5814_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5813_wire_constant, tmp_var);
      BITSEL_u8_u1_5814_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_5824_inst flow-through 
    process(BITSEL_u8_u1_5824_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_5824_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_5823_wire_constant = "& Convert_SLV_To_Hex_String(konst_5823_wire_constant) & " outputs:" & " BITSEL_u8_u1_5824_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_5824_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_5824_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5823_wire_constant, tmp_var);
      BITSEL_u8_u1_5824_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_5834_inst flow-through 
    process(BITSEL_u8_u1_5834_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_5834_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_5833_wire_constant = "& Convert_SLV_To_Hex_String(konst_5833_wire_constant) & " outputs:" & " BITSEL_u8_u1_5834_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_5834_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_5834_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5833_wire_constant, tmp_var);
      BITSEL_u8_u1_5834_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_5844_inst flow-through 
    process(BITSEL_u8_u1_5844_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_5844_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_5843_wire_constant = "& Convert_SLV_To_Hex_String(konst_5843_wire_constant) & " outputs:" & " BITSEL_u8_u1_5844_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_5844_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_5844_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5843_wire_constant, tmp_var);
      BITSEL_u8_u1_5844_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_5854_inst flow-through 
    process(BITSEL_u8_u1_5854_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_5854_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_5853_wire_constant = "& Convert_SLV_To_Hex_String(konst_5853_wire_constant) & " outputs:" & " BITSEL_u8_u1_5854_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_5854_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_5854_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5853_wire_constant, tmp_var);
      BITSEL_u8_u1_5854_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_5864_inst flow-through 
    process(BITSEL_u8_u1_5864_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_5864_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_5863_wire_constant = "& Convert_SLV_To_Hex_String(konst_5863_wire_constant) & " outputs:" & " BITSEL_u8_u1_5864_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_5864_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_5864_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5863_wire_constant, tmp_var);
      BITSEL_u8_u1_5864_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_5874_inst flow-through 
    process(BITSEL_u8_u1_5874_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_5874_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_5873_wire_constant = "& Convert_SLV_To_Hex_String(konst_5873_wire_constant) & " outputs:" & " BITSEL_u8_u1_5874_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_5874_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_5874_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5873_wire_constant, tmp_var);
      BITSEL_u8_u1_5874_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_5884_inst flow-through 
    process(BITSEL_u8_u1_5884_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_5884_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_5883_wire_constant = "& Convert_SLV_To_Hex_String(konst_5883_wire_constant) & " outputs:" & " BITSEL_u8_u1_5884_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_5884_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_5884_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5883_wire_constant, tmp_var);
      BITSEL_u8_u1_5884_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_5894_inst flow-through 
    process(BITSEL_u8_u1_5894_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_5894_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_5893_wire_constant = "& Convert_SLV_To_Hex_String(konst_5893_wire_constant) & " outputs:" & " BITSEL_u8_u1_5894_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_5894_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_5894_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5893_wire_constant, tmp_var);
      BITSEL_u8_u1_5894_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_5902_inst flow-through 
    process(BITSEL_u8_u1_5902_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_5902_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_5901_wire_constant = "& Convert_SLV_To_Hex_String(konst_5901_wire_constant) & " outputs:" & " BITSEL_u8_u1_5902_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_5902_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_5902_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5901_wire_constant, tmp_var);
      BITSEL_u8_u1_5902_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_5910_inst flow-through 
    process(BITSEL_u8_u1_5910_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_5910_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_5909_wire_constant = "& Convert_SLV_To_Hex_String(konst_5909_wire_constant) & " outputs:" & " BITSEL_u8_u1_5910_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_5910_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_5910_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5909_wire_constant, tmp_var);
      BITSEL_u8_u1_5910_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_5918_inst flow-through 
    process(BITSEL_u8_u1_5918_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_5918_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_5917_wire_constant = "& Convert_SLV_To_Hex_String(konst_5917_wire_constant) & " outputs:" & " BITSEL_u8_u1_5918_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_5918_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_5918_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5917_wire_constant, tmp_var);
      BITSEL_u8_u1_5918_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_5926_inst flow-through 
    process(BITSEL_u8_u1_5926_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_5926_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_5925_wire_constant = "& Convert_SLV_To_Hex_String(konst_5925_wire_constant) & " outputs:" & " BITSEL_u8_u1_5926_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_5926_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_5926_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5925_wire_constant, tmp_var);
      BITSEL_u8_u1_5926_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_5934_inst flow-through 
    process(BITSEL_u8_u1_5934_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_5934_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_5933_wire_constant = "& Convert_SLV_To_Hex_String(konst_5933_wire_constant) & " outputs:" & " BITSEL_u8_u1_5934_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_5934_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_5934_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5933_wire_constant, tmp_var);
      BITSEL_u8_u1_5934_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_5942_inst flow-through 
    process(BITSEL_u8_u1_5942_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_5942_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_5941_wire_constant = "& Convert_SLV_To_Hex_String(konst_5941_wire_constant) & " outputs:" & " BITSEL_u8_u1_5942_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_5942_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_5942_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5941_wire_constant, tmp_var);
      BITSEL_u8_u1_5942_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_5950_inst flow-through 
    process(BITSEL_u8_u1_5950_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_5950_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_5949_wire_constant = "& Convert_SLV_To_Hex_String(konst_5949_wire_constant) & " outputs:" & " BITSEL_u8_u1_5950_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_5950_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_5950_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5949_wire_constant, tmp_var);
      BITSEL_u8_u1_5950_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_5958_inst flow-through 
    process(BITSEL_u8_u1_5958_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_5958_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_5957_wire_constant = "& Convert_SLV_To_Hex_String(konst_5957_wire_constant) & " outputs:" & " BITSEL_u8_u1_5958_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_5958_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_5958_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5957_wire_constant, tmp_var);
      BITSEL_u8_u1_5958_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_5966_inst flow-through 
    process(BITSEL_u8_u1_5966_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_5966_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_5965_wire_constant = "& Convert_SLV_To_Hex_String(konst_5965_wire_constant) & " outputs:" & " BITSEL_u8_u1_5966_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_5966_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_5966_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5965_wire_constant, tmp_var);
      BITSEL_u8_u1_5966_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_5974_inst flow-through 
    process(BITSEL_u8_u1_5974_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_5974_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_5973_wire_constant = "& Convert_SLV_To_Hex_String(konst_5973_wire_constant) & " outputs:" & " BITSEL_u8_u1_5974_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_5974_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_5974_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5973_wire_constant, tmp_var);
      BITSEL_u8_u1_5974_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_5982_inst flow-through 
    process(BITSEL_u8_u1_5982_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_5982_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_5981_wire_constant = "& Convert_SLV_To_Hex_String(konst_5981_wire_constant) & " outputs:" & " BITSEL_u8_u1_5982_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_5982_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_5982_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5981_wire_constant, tmp_var);
      BITSEL_u8_u1_5982_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_5990_inst flow-through 
    process(BITSEL_u8_u1_5990_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_5990_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_5989_wire_constant = "& Convert_SLV_To_Hex_String(konst_5989_wire_constant) & " outputs:" & " BITSEL_u8_u1_5990_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_5990_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_5990_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5989_wire_constant, tmp_var);
      BITSEL_u8_u1_5990_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_5998_inst flow-through 
    process(BITSEL_u8_u1_5998_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_5998_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_5997_wire_constant = "& Convert_SLV_To_Hex_String(konst_5997_wire_constant) & " outputs:" & " BITSEL_u8_u1_5998_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_5998_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_5998_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5997_wire_constant, tmp_var);
      BITSEL_u8_u1_5998_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6006_inst flow-through 
    process(BITSEL_u8_u1_6006_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6006_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6005_wire_constant = "& Convert_SLV_To_Hex_String(konst_6005_wire_constant) & " outputs:" & " BITSEL_u8_u1_6006_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6006_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6006_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6005_wire_constant, tmp_var);
      BITSEL_u8_u1_6006_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6014_inst flow-through 
    process(BITSEL_u8_u1_6014_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6014_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6013_wire_constant = "& Convert_SLV_To_Hex_String(konst_6013_wire_constant) & " outputs:" & " BITSEL_u8_u1_6014_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6014_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6014_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6013_wire_constant, tmp_var);
      BITSEL_u8_u1_6014_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6022_inst flow-through 
    process(BITSEL_u8_u1_6022_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6022_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6021_wire_constant = "& Convert_SLV_To_Hex_String(konst_6021_wire_constant) & " outputs:" & " BITSEL_u8_u1_6022_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6022_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6022_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6021_wire_constant, tmp_var);
      BITSEL_u8_u1_6022_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6030_inst flow-through 
    process(BITSEL_u8_u1_6030_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6030_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6029_wire_constant = "& Convert_SLV_To_Hex_String(konst_6029_wire_constant) & " outputs:" & " BITSEL_u8_u1_6030_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6030_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6030_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6029_wire_constant, tmp_var);
      BITSEL_u8_u1_6030_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6038_inst flow-through 
    process(BITSEL_u8_u1_6038_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6038_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6037_wire_constant = "& Convert_SLV_To_Hex_String(konst_6037_wire_constant) & " outputs:" & " BITSEL_u8_u1_6038_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6038_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6038_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6037_wire_constant, tmp_var);
      BITSEL_u8_u1_6038_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6046_inst flow-through 
    process(BITSEL_u8_u1_6046_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6046_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6045_wire_constant = "& Convert_SLV_To_Hex_String(konst_6045_wire_constant) & " outputs:" & " BITSEL_u8_u1_6046_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6046_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6046_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6045_wire_constant, tmp_var);
      BITSEL_u8_u1_6046_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6054_inst flow-through 
    process(BITSEL_u8_u1_6054_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6054_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6053_wire_constant = "& Convert_SLV_To_Hex_String(konst_6053_wire_constant) & " outputs:" & " BITSEL_u8_u1_6054_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6054_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6054_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6053_wire_constant, tmp_var);
      BITSEL_u8_u1_6054_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6062_inst flow-through 
    process(BITSEL_u8_u1_6062_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6062_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6061_wire_constant = "& Convert_SLV_To_Hex_String(konst_6061_wire_constant) & " outputs:" & " BITSEL_u8_u1_6062_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6062_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6062_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6061_wire_constant, tmp_var);
      BITSEL_u8_u1_6062_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6070_inst flow-through 
    process(BITSEL_u8_u1_6070_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6070_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6069_wire_constant = "& Convert_SLV_To_Hex_String(konst_6069_wire_constant) & " outputs:" & " BITSEL_u8_u1_6070_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6070_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6070_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6069_wire_constant, tmp_var);
      BITSEL_u8_u1_6070_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6078_inst flow-through 
    process(BITSEL_u8_u1_6078_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6078_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6077_wire_constant = "& Convert_SLV_To_Hex_String(konst_6077_wire_constant) & " outputs:" & " BITSEL_u8_u1_6078_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6078_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6078_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6077_wire_constant, tmp_var);
      BITSEL_u8_u1_6078_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6086_inst flow-through 
    process(BITSEL_u8_u1_6086_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6086_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6085_wire_constant = "& Convert_SLV_To_Hex_String(konst_6085_wire_constant) & " outputs:" & " BITSEL_u8_u1_6086_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6086_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6086_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6085_wire_constant, tmp_var);
      BITSEL_u8_u1_6086_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6094_inst flow-through 
    process(BITSEL_u8_u1_6094_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6094_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6093_wire_constant = "& Convert_SLV_To_Hex_String(konst_6093_wire_constant) & " outputs:" & " BITSEL_u8_u1_6094_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6094_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6094_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6093_wire_constant, tmp_var);
      BITSEL_u8_u1_6094_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6102_inst flow-through 
    process(BITSEL_u8_u1_6102_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6102_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6101_wire_constant = "& Convert_SLV_To_Hex_String(konst_6101_wire_constant) & " outputs:" & " BITSEL_u8_u1_6102_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6102_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6102_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6101_wire_constant, tmp_var);
      BITSEL_u8_u1_6102_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6110_inst flow-through 
    process(BITSEL_u8_u1_6110_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6110_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6109_wire_constant = "& Convert_SLV_To_Hex_String(konst_6109_wire_constant) & " outputs:" & " BITSEL_u8_u1_6110_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6110_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6110_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6109_wire_constant, tmp_var);
      BITSEL_u8_u1_6110_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6118_inst flow-through 
    process(BITSEL_u8_u1_6118_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6118_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6117_wire_constant = "& Convert_SLV_To_Hex_String(konst_6117_wire_constant) & " outputs:" & " BITSEL_u8_u1_6118_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6118_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6118_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6117_wire_constant, tmp_var);
      BITSEL_u8_u1_6118_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6126_inst flow-through 
    process(BITSEL_u8_u1_6126_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6126_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6125_wire_constant = "& Convert_SLV_To_Hex_String(konst_6125_wire_constant) & " outputs:" & " BITSEL_u8_u1_6126_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6126_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6126_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6125_wire_constant, tmp_var);
      BITSEL_u8_u1_6126_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6134_inst flow-through 
    process(BITSEL_u8_u1_6134_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6134_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6133_wire_constant = "& Convert_SLV_To_Hex_String(konst_6133_wire_constant) & " outputs:" & " BITSEL_u8_u1_6134_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6134_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6134_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6133_wire_constant, tmp_var);
      BITSEL_u8_u1_6134_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6142_inst flow-through 
    process(BITSEL_u8_u1_6142_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6142_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6141_wire_constant = "& Convert_SLV_To_Hex_String(konst_6141_wire_constant) & " outputs:" & " BITSEL_u8_u1_6142_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6142_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6142_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6141_wire_constant, tmp_var);
      BITSEL_u8_u1_6142_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6150_inst flow-through 
    process(BITSEL_u8_u1_6150_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6150_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6149_wire_constant = "& Convert_SLV_To_Hex_String(konst_6149_wire_constant) & " outputs:" & " BITSEL_u8_u1_6150_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6150_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6150_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6149_wire_constant, tmp_var);
      BITSEL_u8_u1_6150_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6158_inst flow-through 
    process(BITSEL_u8_u1_6158_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6158_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6157_wire_constant = "& Convert_SLV_To_Hex_String(konst_6157_wire_constant) & " outputs:" & " BITSEL_u8_u1_6158_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6158_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6158_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6157_wire_constant, tmp_var);
      BITSEL_u8_u1_6158_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6166_inst flow-through 
    process(BITSEL_u8_u1_6166_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6166_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6165_wire_constant = "& Convert_SLV_To_Hex_String(konst_6165_wire_constant) & " outputs:" & " BITSEL_u8_u1_6166_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6166_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6166_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6165_wire_constant, tmp_var);
      BITSEL_u8_u1_6166_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6174_inst flow-through 
    process(BITSEL_u8_u1_6174_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6174_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6173_wire_constant = "& Convert_SLV_To_Hex_String(konst_6173_wire_constant) & " outputs:" & " BITSEL_u8_u1_6174_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6174_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6174_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6173_wire_constant, tmp_var);
      BITSEL_u8_u1_6174_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6182_inst flow-through 
    process(BITSEL_u8_u1_6182_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6182_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6181_wire_constant = "& Convert_SLV_To_Hex_String(konst_6181_wire_constant) & " outputs:" & " BITSEL_u8_u1_6182_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6182_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6182_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6181_wire_constant, tmp_var);
      BITSEL_u8_u1_6182_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6190_inst flow-through 
    process(BITSEL_u8_u1_6190_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6190_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6189_wire_constant = "& Convert_SLV_To_Hex_String(konst_6189_wire_constant) & " outputs:" & " BITSEL_u8_u1_6190_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6190_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6190_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6189_wire_constant, tmp_var);
      BITSEL_u8_u1_6190_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6198_inst flow-through 
    process(BITSEL_u8_u1_6198_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6198_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6197_wire_constant = "& Convert_SLV_To_Hex_String(konst_6197_wire_constant) & " outputs:" & " BITSEL_u8_u1_6198_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6198_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6198_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6197_wire_constant, tmp_var);
      BITSEL_u8_u1_6198_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6206_inst flow-through 
    process(BITSEL_u8_u1_6206_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6206_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6205_wire_constant = "& Convert_SLV_To_Hex_String(konst_6205_wire_constant) & " outputs:" & " BITSEL_u8_u1_6206_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6206_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6206_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6205_wire_constant, tmp_var);
      BITSEL_u8_u1_6206_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6214_inst flow-through 
    process(BITSEL_u8_u1_6214_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6214_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6213_wire_constant = "& Convert_SLV_To_Hex_String(konst_6213_wire_constant) & " outputs:" & " BITSEL_u8_u1_6214_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6214_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6214_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6213_wire_constant, tmp_var);
      BITSEL_u8_u1_6214_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6222_inst flow-through 
    process(BITSEL_u8_u1_6222_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6222_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6221_wire_constant = "& Convert_SLV_To_Hex_String(konst_6221_wire_constant) & " outputs:" & " BITSEL_u8_u1_6222_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6222_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6222_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6221_wire_constant, tmp_var);
      BITSEL_u8_u1_6222_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6230_inst flow-through 
    process(BITSEL_u8_u1_6230_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6230_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6229_wire_constant = "& Convert_SLV_To_Hex_String(konst_6229_wire_constant) & " outputs:" & " BITSEL_u8_u1_6230_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6230_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6230_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6229_wire_constant, tmp_var);
      BITSEL_u8_u1_6230_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6238_inst flow-through 
    process(BITSEL_u8_u1_6238_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6238_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6237_wire_constant = "& Convert_SLV_To_Hex_String(konst_6237_wire_constant) & " outputs:" & " BITSEL_u8_u1_6238_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6238_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6238_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6237_wire_constant, tmp_var);
      BITSEL_u8_u1_6238_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6246_inst flow-through 
    process(BITSEL_u8_u1_6246_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6246_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6245_wire_constant = "& Convert_SLV_To_Hex_String(konst_6245_wire_constant) & " outputs:" & " BITSEL_u8_u1_6246_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6246_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6246_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6245_wire_constant, tmp_var);
      BITSEL_u8_u1_6246_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6254_inst flow-through 
    process(BITSEL_u8_u1_6254_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6254_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6253_wire_constant = "& Convert_SLV_To_Hex_String(konst_6253_wire_constant) & " outputs:" & " BITSEL_u8_u1_6254_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6254_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6254_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6253_wire_constant, tmp_var);
      BITSEL_u8_u1_6254_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6262_inst flow-through 
    process(BITSEL_u8_u1_6262_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6262_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6261_wire_constant = "& Convert_SLV_To_Hex_String(konst_6261_wire_constant) & " outputs:" & " BITSEL_u8_u1_6262_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6262_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6262_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6261_wire_constant, tmp_var);
      BITSEL_u8_u1_6262_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6270_inst flow-through 
    process(BITSEL_u8_u1_6270_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6270_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6269_wire_constant = "& Convert_SLV_To_Hex_String(konst_6269_wire_constant) & " outputs:" & " BITSEL_u8_u1_6270_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6270_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6270_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6269_wire_constant, tmp_var);
      BITSEL_u8_u1_6270_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6278_inst flow-through 
    process(BITSEL_u8_u1_6278_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6278_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6277_wire_constant = "& Convert_SLV_To_Hex_String(konst_6277_wire_constant) & " outputs:" & " BITSEL_u8_u1_6278_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6278_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6278_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6277_wire_constant, tmp_var);
      BITSEL_u8_u1_6278_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6286_inst flow-through 
    process(BITSEL_u8_u1_6286_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6286_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6285_wire_constant = "& Convert_SLV_To_Hex_String(konst_6285_wire_constant) & " outputs:" & " BITSEL_u8_u1_6286_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6286_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6286_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6285_wire_constant, tmp_var);
      BITSEL_u8_u1_6286_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6294_inst flow-through 
    process(BITSEL_u8_u1_6294_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6294_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6293_wire_constant = "& Convert_SLV_To_Hex_String(konst_6293_wire_constant) & " outputs:" & " BITSEL_u8_u1_6294_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6294_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6294_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6293_wire_constant, tmp_var);
      BITSEL_u8_u1_6294_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6302_inst flow-through 
    process(BITSEL_u8_u1_6302_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6302_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6301_wire_constant = "& Convert_SLV_To_Hex_String(konst_6301_wire_constant) & " outputs:" & " BITSEL_u8_u1_6302_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6302_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6302_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6301_wire_constant, tmp_var);
      BITSEL_u8_u1_6302_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6310_inst flow-through 
    process(BITSEL_u8_u1_6310_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6310_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6309_wire_constant = "& Convert_SLV_To_Hex_String(konst_6309_wire_constant) & " outputs:" & " BITSEL_u8_u1_6310_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6310_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6310_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6309_wire_constant, tmp_var);
      BITSEL_u8_u1_6310_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6318_inst flow-through 
    process(BITSEL_u8_u1_6318_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6318_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6317_wire_constant = "& Convert_SLV_To_Hex_String(konst_6317_wire_constant) & " outputs:" & " BITSEL_u8_u1_6318_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6318_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6318_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6317_wire_constant, tmp_var);
      BITSEL_u8_u1_6318_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6326_inst flow-through 
    process(BITSEL_u8_u1_6326_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6326_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6325_wire_constant = "& Convert_SLV_To_Hex_String(konst_6325_wire_constant) & " outputs:" & " BITSEL_u8_u1_6326_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6326_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6326_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6325_wire_constant, tmp_var);
      BITSEL_u8_u1_6326_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6334_inst flow-through 
    process(BITSEL_u8_u1_6334_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6334_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6333_wire_constant = "& Convert_SLV_To_Hex_String(konst_6333_wire_constant) & " outputs:" & " BITSEL_u8_u1_6334_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6334_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6334_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6333_wire_constant, tmp_var);
      BITSEL_u8_u1_6334_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6342_inst flow-through 
    process(BITSEL_u8_u1_6342_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6342_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6341_wire_constant = "& Convert_SLV_To_Hex_String(konst_6341_wire_constant) & " outputs:" & " BITSEL_u8_u1_6342_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6342_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6342_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6341_wire_constant, tmp_var);
      BITSEL_u8_u1_6342_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6350_inst flow-through 
    process(BITSEL_u8_u1_6350_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6350_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6349_wire_constant = "& Convert_SLV_To_Hex_String(konst_6349_wire_constant) & " outputs:" & " BITSEL_u8_u1_6350_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6350_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6350_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6349_wire_constant, tmp_var);
      BITSEL_u8_u1_6350_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6358_inst flow-through 
    process(BITSEL_u8_u1_6358_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6358_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6357_wire_constant = "& Convert_SLV_To_Hex_String(konst_6357_wire_constant) & " outputs:" & " BITSEL_u8_u1_6358_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6358_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6358_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6357_wire_constant, tmp_var);
      BITSEL_u8_u1_6358_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6366_inst flow-through 
    process(BITSEL_u8_u1_6366_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6366_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6365_wire_constant = "& Convert_SLV_To_Hex_String(konst_6365_wire_constant) & " outputs:" & " BITSEL_u8_u1_6366_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6366_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6366_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6365_wire_constant, tmp_var);
      BITSEL_u8_u1_6366_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6374_inst flow-through 
    process(BITSEL_u8_u1_6374_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6374_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6373_wire_constant = "& Convert_SLV_To_Hex_String(konst_6373_wire_constant) & " outputs:" & " BITSEL_u8_u1_6374_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6374_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6374_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6373_wire_constant, tmp_var);
      BITSEL_u8_u1_6374_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6382_inst flow-through 
    process(BITSEL_u8_u1_6382_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6382_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6381_wire_constant = "& Convert_SLV_To_Hex_String(konst_6381_wire_constant) & " outputs:" & " BITSEL_u8_u1_6382_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6382_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6382_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6381_wire_constant, tmp_var);
      BITSEL_u8_u1_6382_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6390_inst flow-through 
    process(BITSEL_u8_u1_6390_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6390_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6389_wire_constant = "& Convert_SLV_To_Hex_String(konst_6389_wire_constant) & " outputs:" & " BITSEL_u8_u1_6390_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6390_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6390_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6389_wire_constant, tmp_var);
      BITSEL_u8_u1_6390_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6398_inst flow-through 
    process(BITSEL_u8_u1_6398_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6398_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6397_wire_constant = "& Convert_SLV_To_Hex_String(konst_6397_wire_constant) & " outputs:" & " BITSEL_u8_u1_6398_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6398_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6398_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6397_wire_constant, tmp_var);
      BITSEL_u8_u1_6398_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6406_inst flow-through 
    process(BITSEL_u8_u1_6406_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6406_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6405_wire_constant = "& Convert_SLV_To_Hex_String(konst_6405_wire_constant) & " outputs:" & " BITSEL_u8_u1_6406_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6406_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6406_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6405_wire_constant, tmp_var);
      BITSEL_u8_u1_6406_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6414_inst flow-through 
    process(BITSEL_u8_u1_6414_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6414_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6413_wire_constant = "& Convert_SLV_To_Hex_String(konst_6413_wire_constant) & " outputs:" & " BITSEL_u8_u1_6414_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6414_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6414_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6413_wire_constant, tmp_var);
      BITSEL_u8_u1_6414_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6422_inst flow-through 
    process(BITSEL_u8_u1_6422_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6422_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6421_wire_constant = "& Convert_SLV_To_Hex_String(konst_6421_wire_constant) & " outputs:" & " BITSEL_u8_u1_6422_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6422_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6422_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6421_wire_constant, tmp_var);
      BITSEL_u8_u1_6422_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6430_inst flow-through 
    process(BITSEL_u8_u1_6430_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6430_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6429_wire_constant = "& Convert_SLV_To_Hex_String(konst_6429_wire_constant) & " outputs:" & " BITSEL_u8_u1_6430_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6430_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6430_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6429_wire_constant, tmp_var);
      BITSEL_u8_u1_6430_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6438_inst flow-through 
    process(BITSEL_u8_u1_6438_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6438_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6437_wire_constant = "& Convert_SLV_To_Hex_String(konst_6437_wire_constant) & " outputs:" & " BITSEL_u8_u1_6438_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6438_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6438_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6437_wire_constant, tmp_var);
      BITSEL_u8_u1_6438_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6446_inst flow-through 
    process(BITSEL_u8_u1_6446_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6446_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6445_wire_constant = "& Convert_SLV_To_Hex_String(konst_6445_wire_constant) & " outputs:" & " BITSEL_u8_u1_6446_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6446_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6446_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6445_wire_constant, tmp_var);
      BITSEL_u8_u1_6446_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6454_inst flow-through 
    process(BITSEL_u8_u1_6454_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6454_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6453_wire_constant = "& Convert_SLV_To_Hex_String(konst_6453_wire_constant) & " outputs:" & " BITSEL_u8_u1_6454_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6454_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6454_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6453_wire_constant, tmp_var);
      BITSEL_u8_u1_6454_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6462_inst flow-through 
    process(BITSEL_u8_u1_6462_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6462_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6461_wire_constant = "& Convert_SLV_To_Hex_String(konst_6461_wire_constant) & " outputs:" & " BITSEL_u8_u1_6462_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6462_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6462_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6461_wire_constant, tmp_var);
      BITSEL_u8_u1_6462_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6470_inst flow-through 
    process(BITSEL_u8_u1_6470_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6470_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6469_wire_constant = "& Convert_SLV_To_Hex_String(konst_6469_wire_constant) & " outputs:" & " BITSEL_u8_u1_6470_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6470_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6470_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6469_wire_constant, tmp_var);
      BITSEL_u8_u1_6470_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6478_inst flow-through 
    process(BITSEL_u8_u1_6478_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6478_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6477_wire_constant = "& Convert_SLV_To_Hex_String(konst_6477_wire_constant) & " outputs:" & " BITSEL_u8_u1_6478_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6478_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6478_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6477_wire_constant, tmp_var);
      BITSEL_u8_u1_6478_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6486_inst flow-through 
    process(BITSEL_u8_u1_6486_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6486_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6485_wire_constant = "& Convert_SLV_To_Hex_String(konst_6485_wire_constant) & " outputs:" & " BITSEL_u8_u1_6486_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6486_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6486_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6485_wire_constant, tmp_var);
      BITSEL_u8_u1_6486_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6494_inst flow-through 
    process(BITSEL_u8_u1_6494_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6494_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6493_wire_constant = "& Convert_SLV_To_Hex_String(konst_6493_wire_constant) & " outputs:" & " BITSEL_u8_u1_6494_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6494_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6494_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6493_wire_constant, tmp_var);
      BITSEL_u8_u1_6494_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6502_inst flow-through 
    process(BITSEL_u8_u1_6502_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6502_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6501_wire_constant = "& Convert_SLV_To_Hex_String(konst_6501_wire_constant) & " outputs:" & " BITSEL_u8_u1_6502_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6502_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6502_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6501_wire_constant, tmp_var);
      BITSEL_u8_u1_6502_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6510_inst flow-through 
    process(BITSEL_u8_u1_6510_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6510_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6509_wire_constant = "& Convert_SLV_To_Hex_String(konst_6509_wire_constant) & " outputs:" & " BITSEL_u8_u1_6510_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6510_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6510_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6509_wire_constant, tmp_var);
      BITSEL_u8_u1_6510_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6518_inst flow-through 
    process(BITSEL_u8_u1_6518_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6518_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6517_wire_constant = "& Convert_SLV_To_Hex_String(konst_6517_wire_constant) & " outputs:" & " BITSEL_u8_u1_6518_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6518_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6518_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6517_wire_constant, tmp_var);
      BITSEL_u8_u1_6518_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6526_inst flow-through 
    process(BITSEL_u8_u1_6526_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6526_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6525_wire_constant = "& Convert_SLV_To_Hex_String(konst_6525_wire_constant) & " outputs:" & " BITSEL_u8_u1_6526_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6526_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6526_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6525_wire_constant, tmp_var);
      BITSEL_u8_u1_6526_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6534_inst flow-through 
    process(BITSEL_u8_u1_6534_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6534_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6533_wire_constant = "& Convert_SLV_To_Hex_String(konst_6533_wire_constant) & " outputs:" & " BITSEL_u8_u1_6534_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6534_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6534_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6533_wire_constant, tmp_var);
      BITSEL_u8_u1_6534_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6542_inst flow-through 
    process(BITSEL_u8_u1_6542_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6542_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6541_wire_constant = "& Convert_SLV_To_Hex_String(konst_6541_wire_constant) & " outputs:" & " BITSEL_u8_u1_6542_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6542_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6542_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6541_wire_constant, tmp_var);
      BITSEL_u8_u1_6542_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6550_inst flow-through 
    process(BITSEL_u8_u1_6550_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6550_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6549_wire_constant = "& Convert_SLV_To_Hex_String(konst_6549_wire_constant) & " outputs:" & " BITSEL_u8_u1_6550_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6550_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6550_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6549_wire_constant, tmp_var);
      BITSEL_u8_u1_6550_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6558_inst flow-through 
    process(BITSEL_u8_u1_6558_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6558_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6557_wire_constant = "& Convert_SLV_To_Hex_String(konst_6557_wire_constant) & " outputs:" & " BITSEL_u8_u1_6558_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6558_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6558_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6557_wire_constant, tmp_var);
      BITSEL_u8_u1_6558_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6566_inst flow-through 
    process(BITSEL_u8_u1_6566_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6566_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6565_wire_constant = "& Convert_SLV_To_Hex_String(konst_6565_wire_constant) & " outputs:" & " BITSEL_u8_u1_6566_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6566_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6566_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6565_wire_constant, tmp_var);
      BITSEL_u8_u1_6566_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6574_inst flow-through 
    process(BITSEL_u8_u1_6574_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6574_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6573_wire_constant = "& Convert_SLV_To_Hex_String(konst_6573_wire_constant) & " outputs:" & " BITSEL_u8_u1_6574_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6574_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6574_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6573_wire_constant, tmp_var);
      BITSEL_u8_u1_6574_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6582_inst flow-through 
    process(BITSEL_u8_u1_6582_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6582_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6581_wire_constant = "& Convert_SLV_To_Hex_String(konst_6581_wire_constant) & " outputs:" & " BITSEL_u8_u1_6582_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6582_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6582_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6581_wire_constant, tmp_var);
      BITSEL_u8_u1_6582_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6590_inst flow-through 
    process(BITSEL_u8_u1_6590_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6590_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6589_wire_constant = "& Convert_SLV_To_Hex_String(konst_6589_wire_constant) & " outputs:" & " BITSEL_u8_u1_6590_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6590_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6590_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6589_wire_constant, tmp_var);
      BITSEL_u8_u1_6590_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6598_inst flow-through 
    process(BITSEL_u8_u1_6598_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6598_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6597_wire_constant = "& Convert_SLV_To_Hex_String(konst_6597_wire_constant) & " outputs:" & " BITSEL_u8_u1_6598_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6598_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6598_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6597_wire_constant, tmp_var);
      BITSEL_u8_u1_6598_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6606_inst flow-through 
    process(BITSEL_u8_u1_6606_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6606_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6605_wire_constant = "& Convert_SLV_To_Hex_String(konst_6605_wire_constant) & " outputs:" & " BITSEL_u8_u1_6606_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6606_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6606_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6605_wire_constant, tmp_var);
      BITSEL_u8_u1_6606_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6614_inst flow-through 
    process(BITSEL_u8_u1_6614_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6614_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6613_wire_constant = "& Convert_SLV_To_Hex_String(konst_6613_wire_constant) & " outputs:" & " BITSEL_u8_u1_6614_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6614_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6614_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6613_wire_constant, tmp_var);
      BITSEL_u8_u1_6614_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6622_inst flow-through 
    process(BITSEL_u8_u1_6622_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6622_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6621_wire_constant = "& Convert_SLV_To_Hex_String(konst_6621_wire_constant) & " outputs:" & " BITSEL_u8_u1_6622_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6622_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6622_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6621_wire_constant, tmp_var);
      BITSEL_u8_u1_6622_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6630_inst flow-through 
    process(BITSEL_u8_u1_6630_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6630_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6629_wire_constant = "& Convert_SLV_To_Hex_String(konst_6629_wire_constant) & " outputs:" & " BITSEL_u8_u1_6630_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6630_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6630_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6629_wire_constant, tmp_var);
      BITSEL_u8_u1_6630_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6638_inst flow-through 
    process(BITSEL_u8_u1_6638_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6638_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6637_wire_constant = "& Convert_SLV_To_Hex_String(konst_6637_wire_constant) & " outputs:" & " BITSEL_u8_u1_6638_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6638_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6638_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6637_wire_constant, tmp_var);
      BITSEL_u8_u1_6638_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6646_inst flow-through 
    process(BITSEL_u8_u1_6646_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6646_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6645_wire_constant = "& Convert_SLV_To_Hex_String(konst_6645_wire_constant) & " outputs:" & " BITSEL_u8_u1_6646_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6646_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6646_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6645_wire_constant, tmp_var);
      BITSEL_u8_u1_6646_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6654_inst flow-through 
    process(BITSEL_u8_u1_6654_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6654_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6653_wire_constant = "& Convert_SLV_To_Hex_String(konst_6653_wire_constant) & " outputs:" & " BITSEL_u8_u1_6654_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6654_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6654_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6653_wire_constant, tmp_var);
      BITSEL_u8_u1_6654_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6662_inst flow-through 
    process(BITSEL_u8_u1_6662_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6662_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6661_wire_constant = "& Convert_SLV_To_Hex_String(konst_6661_wire_constant) & " outputs:" & " BITSEL_u8_u1_6662_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6662_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6662_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6661_wire_constant, tmp_var);
      BITSEL_u8_u1_6662_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6670_inst flow-through 
    process(BITSEL_u8_u1_6670_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6670_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6669_wire_constant = "& Convert_SLV_To_Hex_String(konst_6669_wire_constant) & " outputs:" & " BITSEL_u8_u1_6670_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6670_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6670_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6669_wire_constant, tmp_var);
      BITSEL_u8_u1_6670_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6678_inst flow-through 
    process(BITSEL_u8_u1_6678_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6678_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6677_wire_constant = "& Convert_SLV_To_Hex_String(konst_6677_wire_constant) & " outputs:" & " BITSEL_u8_u1_6678_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6678_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6678_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6677_wire_constant, tmp_var);
      BITSEL_u8_u1_6678_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6686_inst flow-through 
    process(BITSEL_u8_u1_6686_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6686_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6685_wire_constant = "& Convert_SLV_To_Hex_String(konst_6685_wire_constant) & " outputs:" & " BITSEL_u8_u1_6686_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6686_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6686_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6685_wire_constant, tmp_var);
      BITSEL_u8_u1_6686_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6694_inst flow-through 
    process(BITSEL_u8_u1_6694_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6694_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6693_wire_constant = "& Convert_SLV_To_Hex_String(konst_6693_wire_constant) & " outputs:" & " BITSEL_u8_u1_6694_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6694_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6694_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6693_wire_constant, tmp_var);
      BITSEL_u8_u1_6694_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6702_inst flow-through 
    process(BITSEL_u8_u1_6702_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6702_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6701_wire_constant = "& Convert_SLV_To_Hex_String(konst_6701_wire_constant) & " outputs:" & " BITSEL_u8_u1_6702_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6702_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6702_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6701_wire_constant, tmp_var);
      BITSEL_u8_u1_6702_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6710_inst flow-through 
    process(BITSEL_u8_u1_6710_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6710_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6709_wire_constant = "& Convert_SLV_To_Hex_String(konst_6709_wire_constant) & " outputs:" & " BITSEL_u8_u1_6710_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6710_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6710_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6709_wire_constant, tmp_var);
      BITSEL_u8_u1_6710_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6718_inst flow-through 
    process(BITSEL_u8_u1_6718_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6718_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6717_wire_constant = "& Convert_SLV_To_Hex_String(konst_6717_wire_constant) & " outputs:" & " BITSEL_u8_u1_6718_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6718_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6718_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6717_wire_constant, tmp_var);
      BITSEL_u8_u1_6718_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6726_inst flow-through 
    process(BITSEL_u8_u1_6726_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6726_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6725_wire_constant = "& Convert_SLV_To_Hex_String(konst_6725_wire_constant) & " outputs:" & " BITSEL_u8_u1_6726_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6726_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6726_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6725_wire_constant, tmp_var);
      BITSEL_u8_u1_6726_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6734_inst flow-through 
    process(BITSEL_u8_u1_6734_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6734_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6733_wire_constant = "& Convert_SLV_To_Hex_String(konst_6733_wire_constant) & " outputs:" & " BITSEL_u8_u1_6734_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6734_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6734_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6733_wire_constant, tmp_var);
      BITSEL_u8_u1_6734_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6742_inst flow-through 
    process(BITSEL_u8_u1_6742_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6742_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6741_wire_constant = "& Convert_SLV_To_Hex_String(konst_6741_wire_constant) & " outputs:" & " BITSEL_u8_u1_6742_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6742_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6742_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6741_wire_constant, tmp_var);
      BITSEL_u8_u1_6742_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6750_inst flow-through 
    process(BITSEL_u8_u1_6750_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6750_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6749_wire_constant = "& Convert_SLV_To_Hex_String(konst_6749_wire_constant) & " outputs:" & " BITSEL_u8_u1_6750_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6750_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6750_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6749_wire_constant, tmp_var);
      BITSEL_u8_u1_6750_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6758_inst flow-through 
    process(BITSEL_u8_u1_6758_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6758_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6757_wire_constant = "& Convert_SLV_To_Hex_String(konst_6757_wire_constant) & " outputs:" & " BITSEL_u8_u1_6758_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6758_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6758_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6757_wire_constant, tmp_var);
      BITSEL_u8_u1_6758_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6766_inst flow-through 
    process(BITSEL_u8_u1_6766_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6766_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6765_wire_constant = "& Convert_SLV_To_Hex_String(konst_6765_wire_constant) & " outputs:" & " BITSEL_u8_u1_6766_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6766_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6766_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6765_wire_constant, tmp_var);
      BITSEL_u8_u1_6766_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6774_inst flow-through 
    process(BITSEL_u8_u1_6774_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6774_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6773_wire_constant = "& Convert_SLV_To_Hex_String(konst_6773_wire_constant) & " outputs:" & " BITSEL_u8_u1_6774_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6774_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6774_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6773_wire_constant, tmp_var);
      BITSEL_u8_u1_6774_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6782_inst flow-through 
    process(BITSEL_u8_u1_6782_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6782_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6781_wire_constant = "& Convert_SLV_To_Hex_String(konst_6781_wire_constant) & " outputs:" & " BITSEL_u8_u1_6782_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6782_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6782_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6781_wire_constant, tmp_var);
      BITSEL_u8_u1_6782_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6790_inst flow-through 
    process(BITSEL_u8_u1_6790_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6790_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6789_wire_constant = "& Convert_SLV_To_Hex_String(konst_6789_wire_constant) & " outputs:" & " BITSEL_u8_u1_6790_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6790_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6790_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6789_wire_constant, tmp_var);
      BITSEL_u8_u1_6790_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6798_inst flow-through 
    process(BITSEL_u8_u1_6798_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6798_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6797_wire_constant = "& Convert_SLV_To_Hex_String(konst_6797_wire_constant) & " outputs:" & " BITSEL_u8_u1_6798_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6798_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6798_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6797_wire_constant, tmp_var);
      BITSEL_u8_u1_6798_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6806_inst flow-through 
    process(BITSEL_u8_u1_6806_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6806_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6805_wire_constant = "& Convert_SLV_To_Hex_String(konst_6805_wire_constant) & " outputs:" & " BITSEL_u8_u1_6806_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6806_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6806_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6805_wire_constant, tmp_var);
      BITSEL_u8_u1_6806_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6814_inst flow-through 
    process(BITSEL_u8_u1_6814_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6814_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6813_wire_constant = "& Convert_SLV_To_Hex_String(konst_6813_wire_constant) & " outputs:" & " BITSEL_u8_u1_6814_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6814_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6814_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6813_wire_constant, tmp_var);
      BITSEL_u8_u1_6814_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6822_inst flow-through 
    process(BITSEL_u8_u1_6822_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6822_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6821_wire_constant = "& Convert_SLV_To_Hex_String(konst_6821_wire_constant) & " outputs:" & " BITSEL_u8_u1_6822_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6822_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6822_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6821_wire_constant, tmp_var);
      BITSEL_u8_u1_6822_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6830_inst flow-through 
    process(BITSEL_u8_u1_6830_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6830_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6829_wire_constant = "& Convert_SLV_To_Hex_String(konst_6829_wire_constant) & " outputs:" & " BITSEL_u8_u1_6830_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6830_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6830_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6829_wire_constant, tmp_var);
      BITSEL_u8_u1_6830_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6838_inst flow-through 
    process(BITSEL_u8_u1_6838_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6838_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6837_wire_constant = "& Convert_SLV_To_Hex_String(konst_6837_wire_constant) & " outputs:" & " BITSEL_u8_u1_6838_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6838_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6838_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6837_wire_constant, tmp_var);
      BITSEL_u8_u1_6838_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6846_inst flow-through 
    process(BITSEL_u8_u1_6846_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6846_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6845_wire_constant = "& Convert_SLV_To_Hex_String(konst_6845_wire_constant) & " outputs:" & " BITSEL_u8_u1_6846_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6846_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6846_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6845_wire_constant, tmp_var);
      BITSEL_u8_u1_6846_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6854_inst flow-through 
    process(BITSEL_u8_u1_6854_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6854_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6853_wire_constant = "& Convert_SLV_To_Hex_String(konst_6853_wire_constant) & " outputs:" & " BITSEL_u8_u1_6854_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6854_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6854_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6853_wire_constant, tmp_var);
      BITSEL_u8_u1_6854_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6862_inst flow-through 
    process(BITSEL_u8_u1_6862_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6862_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6861_wire_constant = "& Convert_SLV_To_Hex_String(konst_6861_wire_constant) & " outputs:" & " BITSEL_u8_u1_6862_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6862_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6862_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6861_wire_constant, tmp_var);
      BITSEL_u8_u1_6862_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6870_inst flow-through 
    process(BITSEL_u8_u1_6870_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6870_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6869_wire_constant = "& Convert_SLV_To_Hex_String(konst_6869_wire_constant) & " outputs:" & " BITSEL_u8_u1_6870_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6870_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6870_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6869_wire_constant, tmp_var);
      BITSEL_u8_u1_6870_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6878_inst flow-through 
    process(BITSEL_u8_u1_6878_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6878_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6877_wire_constant = "& Convert_SLV_To_Hex_String(konst_6877_wire_constant) & " outputs:" & " BITSEL_u8_u1_6878_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6878_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6878_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6877_wire_constant, tmp_var);
      BITSEL_u8_u1_6878_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6886_inst flow-through 
    process(BITSEL_u8_u1_6886_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6886_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6885_wire_constant = "& Convert_SLV_To_Hex_String(konst_6885_wire_constant) & " outputs:" & " BITSEL_u8_u1_6886_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6886_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6886_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6885_wire_constant, tmp_var);
      BITSEL_u8_u1_6886_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6894_inst flow-through 
    process(BITSEL_u8_u1_6894_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6894_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6893_wire_constant = "& Convert_SLV_To_Hex_String(konst_6893_wire_constant) & " outputs:" & " BITSEL_u8_u1_6894_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6894_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6894_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6893_wire_constant, tmp_var);
      BITSEL_u8_u1_6894_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6902_inst flow-through 
    process(BITSEL_u8_u1_6902_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_3:DP:BITSEL_u8_u1_6902_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6901_wire_constant = "& Convert_SLV_To_Hex_String(konst_6901_wire_constant) & " outputs:" & " BITSEL_u8_u1_6902_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6902_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6902_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6901_wire_constant, tmp_var);
      BITSEL_u8_u1_6902_wire <= tmp_var; -- 
    end process;
    -- 
  end Block; -- data_path
  -- 
end Inv_Sbox_3_Volatile_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library GhdlLink;
use GhdlLink.LogUtilities.all;
library work;
use work.ahir_system_global_package.all;
entity Inv_Sbox_4_Volatile is -- 
  port ( -- 
    clk, reset: in std_logic; 
    s_in : in  std_logic_vector(7 downto 0);
    s_out : out  std_logic_vector(7 downto 0)-- 
  );
  -- 
end entity Inv_Sbox_4_Volatile;
architecture Inv_Sbox_4_Volatile_arch of Inv_Sbox_4_Volatile is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector(8-1 downto 0);
  signal default_zero_sig: std_logic;
  -- input port buffer signals
  signal s_in_buffer :  std_logic_vector(7 downto 0);
  -- output port buffer signals
  signal s_out_buffer :  std_logic_vector(7 downto 0);
  -- volatile/operator module components. 
  signal global_clock_cycle_count: integer := 0;
  -- 
begin --  
  ---------------------------------------------------------- 
  process(clk)  
  begin -- 
    if(clk'event and clk = '1') then -- 
      if(reset = '1') then -- 
        global_clock_cycle_count <= 0; --
      else -- 
        global_clock_cycle_count <= global_clock_cycle_count + 1; -- 
      end if; --
    end if; --
  end process;
  ---------------------------------------------------------- 
  -- input handling ------------------------------------------------
  s_in_buffer <= s_in;
  -- output handling  -------------------------------------------------------
  s_out <= s_out_buffer;
  -- the control path --------------------------------------------------
  default_zero_sig <= '0';
  -- volatile module, no control path
  -- the data path
  data_path: Block -- 
    signal BITSEL_u8_u1_6914_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6924_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6934_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6944_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6954_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6964_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6974_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6984_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6994_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7004_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7014_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7024_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7034_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7044_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7054_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7064_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7074_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7084_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7094_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7104_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7114_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7124_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7134_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7144_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7154_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7164_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7174_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7184_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7194_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7204_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7214_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7224_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7234_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7244_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7254_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7264_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7274_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7284_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7294_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7304_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7314_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7324_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7334_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7344_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7354_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7364_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7374_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7384_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7394_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7404_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7414_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7424_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7434_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7444_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7454_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7464_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7474_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7484_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7494_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7504_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7514_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7524_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7534_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7544_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7554_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7564_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7574_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7584_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7594_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7604_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7614_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7624_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7634_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7644_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7654_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7664_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7674_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7684_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7694_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7704_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7714_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7724_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7734_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7744_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7754_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7764_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7774_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7784_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7794_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7804_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7814_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7824_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7834_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7844_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7854_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7864_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7874_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7884_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7894_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7904_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7914_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7924_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7934_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7944_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7954_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7964_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7974_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7984_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7994_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8004_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8014_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8024_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8034_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8044_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8054_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8064_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8074_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8084_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8094_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8104_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8114_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8124_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8134_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8144_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8154_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8164_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8174_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8184_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8194_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8202_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8210_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8218_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8226_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8234_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8242_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8250_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8258_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8266_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8274_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8282_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8290_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8298_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8306_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8314_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8322_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8330_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8338_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8346_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8354_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8362_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8370_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8378_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8386_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8394_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8402_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8410_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8418_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8426_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8434_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8442_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8450_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8458_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8466_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8474_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8482_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8490_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8498_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8506_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8514_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8522_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8530_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8538_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8546_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8554_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8562_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8570_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8578_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8586_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8594_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8602_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8610_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8618_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8626_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8634_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8642_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8650_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8658_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8666_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8674_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8682_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8690_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8698_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8706_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8714_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8722_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8730_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8738_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8746_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8754_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8762_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8770_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8778_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8786_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8794_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8802_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8810_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8818_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8826_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8834_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8842_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8850_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8858_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8866_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8874_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8882_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8890_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8898_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8906_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8914_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8922_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8930_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8938_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8946_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8954_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8962_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8970_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8978_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8986_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8994_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9002_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9010_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9018_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9026_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9034_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9042_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9050_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9058_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9066_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9074_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9082_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9090_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9098_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9106_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9114_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9122_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9130_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9138_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9146_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9154_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9162_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9170_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9178_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9186_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9194_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9202_wire : std_logic_vector(0 downto 0);
    signal IMA0_6920 : std_logic_vector(7 downto 0);
    signal IMA100_7920 : std_logic_vector(7 downto 0);
    signal IMA101_7930 : std_logic_vector(7 downto 0);
    signal IMA102_7940 : std_logic_vector(7 downto 0);
    signal IMA103_7950 : std_logic_vector(7 downto 0);
    signal IMA104_7960 : std_logic_vector(7 downto 0);
    signal IMA105_7970 : std_logic_vector(7 downto 0);
    signal IMA106_7980 : std_logic_vector(7 downto 0);
    signal IMA107_7990 : std_logic_vector(7 downto 0);
    signal IMA108_8000 : std_logic_vector(7 downto 0);
    signal IMA109_8010 : std_logic_vector(7 downto 0);
    signal IMA10_7020 : std_logic_vector(7 downto 0);
    signal IMA110_8020 : std_logic_vector(7 downto 0);
    signal IMA111_8030 : std_logic_vector(7 downto 0);
    signal IMA112_8040 : std_logic_vector(7 downto 0);
    signal IMA113_8050 : std_logic_vector(7 downto 0);
    signal IMA114_8060 : std_logic_vector(7 downto 0);
    signal IMA115_8070 : std_logic_vector(7 downto 0);
    signal IMA116_8080 : std_logic_vector(7 downto 0);
    signal IMA117_8090 : std_logic_vector(7 downto 0);
    signal IMA118_8100 : std_logic_vector(7 downto 0);
    signal IMA119_8110 : std_logic_vector(7 downto 0);
    signal IMA11_7030 : std_logic_vector(7 downto 0);
    signal IMA120_8120 : std_logic_vector(7 downto 0);
    signal IMA121_8130 : std_logic_vector(7 downto 0);
    signal IMA122_8140 : std_logic_vector(7 downto 0);
    signal IMA123_8150 : std_logic_vector(7 downto 0);
    signal IMA124_8160 : std_logic_vector(7 downto 0);
    signal IMA125_8170 : std_logic_vector(7 downto 0);
    signal IMA126_8180 : std_logic_vector(7 downto 0);
    signal IMA127_8190 : std_logic_vector(7 downto 0);
    signal IMA12_7040 : std_logic_vector(7 downto 0);
    signal IMA13_7050 : std_logic_vector(7 downto 0);
    signal IMA14_7060 : std_logic_vector(7 downto 0);
    signal IMA15_7070 : std_logic_vector(7 downto 0);
    signal IMA16_7080 : std_logic_vector(7 downto 0);
    signal IMA17_7090 : std_logic_vector(7 downto 0);
    signal IMA18_7100 : std_logic_vector(7 downto 0);
    signal IMA19_7110 : std_logic_vector(7 downto 0);
    signal IMA1_6930 : std_logic_vector(7 downto 0);
    signal IMA20_7120 : std_logic_vector(7 downto 0);
    signal IMA21_7130 : std_logic_vector(7 downto 0);
    signal IMA22_7140 : std_logic_vector(7 downto 0);
    signal IMA23_7150 : std_logic_vector(7 downto 0);
    signal IMA24_7160 : std_logic_vector(7 downto 0);
    signal IMA25_7170 : std_logic_vector(7 downto 0);
    signal IMA26_7180 : std_logic_vector(7 downto 0);
    signal IMA27_7190 : std_logic_vector(7 downto 0);
    signal IMA28_7200 : std_logic_vector(7 downto 0);
    signal IMA29_7210 : std_logic_vector(7 downto 0);
    signal IMA2_6940 : std_logic_vector(7 downto 0);
    signal IMA30_7220 : std_logic_vector(7 downto 0);
    signal IMA31_7230 : std_logic_vector(7 downto 0);
    signal IMA32_7240 : std_logic_vector(7 downto 0);
    signal IMA33_7250 : std_logic_vector(7 downto 0);
    signal IMA34_7260 : std_logic_vector(7 downto 0);
    signal IMA35_7270 : std_logic_vector(7 downto 0);
    signal IMA36_7280 : std_logic_vector(7 downto 0);
    signal IMA37_7290 : std_logic_vector(7 downto 0);
    signal IMA38_7300 : std_logic_vector(7 downto 0);
    signal IMA39_7310 : std_logic_vector(7 downto 0);
    signal IMA3_6950 : std_logic_vector(7 downto 0);
    signal IMA40_7320 : std_logic_vector(7 downto 0);
    signal IMA41_7330 : std_logic_vector(7 downto 0);
    signal IMA42_7340 : std_logic_vector(7 downto 0);
    signal IMA43_7350 : std_logic_vector(7 downto 0);
    signal IMA44_7360 : std_logic_vector(7 downto 0);
    signal IMA45_7370 : std_logic_vector(7 downto 0);
    signal IMA46_7380 : std_logic_vector(7 downto 0);
    signal IMA47_7390 : std_logic_vector(7 downto 0);
    signal IMA48_7400 : std_logic_vector(7 downto 0);
    signal IMA49_7410 : std_logic_vector(7 downto 0);
    signal IMA4_6960 : std_logic_vector(7 downto 0);
    signal IMA50_7420 : std_logic_vector(7 downto 0);
    signal IMA51_7430 : std_logic_vector(7 downto 0);
    signal IMA52_7440 : std_logic_vector(7 downto 0);
    signal IMA53_7450 : std_logic_vector(7 downto 0);
    signal IMA54_7460 : std_logic_vector(7 downto 0);
    signal IMA55_7470 : std_logic_vector(7 downto 0);
    signal IMA56_7480 : std_logic_vector(7 downto 0);
    signal IMA57_7490 : std_logic_vector(7 downto 0);
    signal IMA58_7500 : std_logic_vector(7 downto 0);
    signal IMA59_7510 : std_logic_vector(7 downto 0);
    signal IMA5_6970 : std_logic_vector(7 downto 0);
    signal IMA60_7520 : std_logic_vector(7 downto 0);
    signal IMA61_7530 : std_logic_vector(7 downto 0);
    signal IMA62_7540 : std_logic_vector(7 downto 0);
    signal IMA63_7550 : std_logic_vector(7 downto 0);
    signal IMA64_7560 : std_logic_vector(7 downto 0);
    signal IMA65_7570 : std_logic_vector(7 downto 0);
    signal IMA66_7580 : std_logic_vector(7 downto 0);
    signal IMA67_7590 : std_logic_vector(7 downto 0);
    signal IMA68_7600 : std_logic_vector(7 downto 0);
    signal IMA69_7610 : std_logic_vector(7 downto 0);
    signal IMA6_6980 : std_logic_vector(7 downto 0);
    signal IMA70_7620 : std_logic_vector(7 downto 0);
    signal IMA71_7630 : std_logic_vector(7 downto 0);
    signal IMA72_7640 : std_logic_vector(7 downto 0);
    signal IMA73_7650 : std_logic_vector(7 downto 0);
    signal IMA74_7660 : std_logic_vector(7 downto 0);
    signal IMA75_7670 : std_logic_vector(7 downto 0);
    signal IMA76_7680 : std_logic_vector(7 downto 0);
    signal IMA77_7690 : std_logic_vector(7 downto 0);
    signal IMA78_7700 : std_logic_vector(7 downto 0);
    signal IMA79_7710 : std_logic_vector(7 downto 0);
    signal IMA7_6990 : std_logic_vector(7 downto 0);
    signal IMA80_7720 : std_logic_vector(7 downto 0);
    signal IMA81_7730 : std_logic_vector(7 downto 0);
    signal IMA82_7740 : std_logic_vector(7 downto 0);
    signal IMA83_7750 : std_logic_vector(7 downto 0);
    signal IMA84_7760 : std_logic_vector(7 downto 0);
    signal IMA85_7770 : std_logic_vector(7 downto 0);
    signal IMA86_7780 : std_logic_vector(7 downto 0);
    signal IMA87_7790 : std_logic_vector(7 downto 0);
    signal IMA88_7800 : std_logic_vector(7 downto 0);
    signal IMA89_7810 : std_logic_vector(7 downto 0);
    signal IMA8_7000 : std_logic_vector(7 downto 0);
    signal IMA90_7820 : std_logic_vector(7 downto 0);
    signal IMA91_7830 : std_logic_vector(7 downto 0);
    signal IMA92_7840 : std_logic_vector(7 downto 0);
    signal IMA93_7850 : std_logic_vector(7 downto 0);
    signal IMA94_7860 : std_logic_vector(7 downto 0);
    signal IMA95_7870 : std_logic_vector(7 downto 0);
    signal IMA96_7880 : std_logic_vector(7 downto 0);
    signal IMA97_7890 : std_logic_vector(7 downto 0);
    signal IMA98_7900 : std_logic_vector(7 downto 0);
    signal IMA99_7910 : std_logic_vector(7 downto 0);
    signal IMA9_7010 : std_logic_vector(7 downto 0);
    signal IMB0_8198 : std_logic_vector(7 downto 0);
    signal IMB10_8278 : std_logic_vector(7 downto 0);
    signal IMB11_8286 : std_logic_vector(7 downto 0);
    signal IMB12_8294 : std_logic_vector(7 downto 0);
    signal IMB13_8302 : std_logic_vector(7 downto 0);
    signal IMB14_8310 : std_logic_vector(7 downto 0);
    signal IMB15_8318 : std_logic_vector(7 downto 0);
    signal IMB16_8326 : std_logic_vector(7 downto 0);
    signal IMB17_8334 : std_logic_vector(7 downto 0);
    signal IMB18_8342 : std_logic_vector(7 downto 0);
    signal IMB19_8350 : std_logic_vector(7 downto 0);
    signal IMB1_8206 : std_logic_vector(7 downto 0);
    signal IMB20_8358 : std_logic_vector(7 downto 0);
    signal IMB21_8366 : std_logic_vector(7 downto 0);
    signal IMB22_8374 : std_logic_vector(7 downto 0);
    signal IMB23_8382 : std_logic_vector(7 downto 0);
    signal IMB24_8390 : std_logic_vector(7 downto 0);
    signal IMB25_8398 : std_logic_vector(7 downto 0);
    signal IMB26_8406 : std_logic_vector(7 downto 0);
    signal IMB27_8414 : std_logic_vector(7 downto 0);
    signal IMB28_8422 : std_logic_vector(7 downto 0);
    signal IMB29_8430 : std_logic_vector(7 downto 0);
    signal IMB2_8214 : std_logic_vector(7 downto 0);
    signal IMB30_8438 : std_logic_vector(7 downto 0);
    signal IMB31_8446 : std_logic_vector(7 downto 0);
    signal IMB32_8454 : std_logic_vector(7 downto 0);
    signal IMB33_8462 : std_logic_vector(7 downto 0);
    signal IMB34_8470 : std_logic_vector(7 downto 0);
    signal IMB35_8478 : std_logic_vector(7 downto 0);
    signal IMB36_8486 : std_logic_vector(7 downto 0);
    signal IMB37_8494 : std_logic_vector(7 downto 0);
    signal IMB38_8502 : std_logic_vector(7 downto 0);
    signal IMB39_8510 : std_logic_vector(7 downto 0);
    signal IMB3_8222 : std_logic_vector(7 downto 0);
    signal IMB40_8518 : std_logic_vector(7 downto 0);
    signal IMB41_8526 : std_logic_vector(7 downto 0);
    signal IMB42_8534 : std_logic_vector(7 downto 0);
    signal IMB43_8542 : std_logic_vector(7 downto 0);
    signal IMB44_8550 : std_logic_vector(7 downto 0);
    signal IMB45_8558 : std_logic_vector(7 downto 0);
    signal IMB46_8566 : std_logic_vector(7 downto 0);
    signal IMB47_8574 : std_logic_vector(7 downto 0);
    signal IMB48_8582 : std_logic_vector(7 downto 0);
    signal IMB49_8590 : std_logic_vector(7 downto 0);
    signal IMB4_8230 : std_logic_vector(7 downto 0);
    signal IMB50_8598 : std_logic_vector(7 downto 0);
    signal IMB51_8606 : std_logic_vector(7 downto 0);
    signal IMB52_8614 : std_logic_vector(7 downto 0);
    signal IMB53_8622 : std_logic_vector(7 downto 0);
    signal IMB54_8630 : std_logic_vector(7 downto 0);
    signal IMB55_8638 : std_logic_vector(7 downto 0);
    signal IMB56_8646 : std_logic_vector(7 downto 0);
    signal IMB57_8654 : std_logic_vector(7 downto 0);
    signal IMB58_8662 : std_logic_vector(7 downto 0);
    signal IMB59_8670 : std_logic_vector(7 downto 0);
    signal IMB5_8238 : std_logic_vector(7 downto 0);
    signal IMB60_8678 : std_logic_vector(7 downto 0);
    signal IMB61_8686 : std_logic_vector(7 downto 0);
    signal IMB62_8694 : std_logic_vector(7 downto 0);
    signal IMB63_8702 : std_logic_vector(7 downto 0);
    signal IMB6_8246 : std_logic_vector(7 downto 0);
    signal IMB7_8254 : std_logic_vector(7 downto 0);
    signal IMB8_8262 : std_logic_vector(7 downto 0);
    signal IMB9_8270 : std_logic_vector(7 downto 0);
    signal IMC0_8710 : std_logic_vector(7 downto 0);
    signal IMC10_8790 : std_logic_vector(7 downto 0);
    signal IMC11_8798 : std_logic_vector(7 downto 0);
    signal IMC12_8806 : std_logic_vector(7 downto 0);
    signal IMC13_8814 : std_logic_vector(7 downto 0);
    signal IMC14_8822 : std_logic_vector(7 downto 0);
    signal IMC15_8830 : std_logic_vector(7 downto 0);
    signal IMC16_8838 : std_logic_vector(7 downto 0);
    signal IMC17_8846 : std_logic_vector(7 downto 0);
    signal IMC18_8854 : std_logic_vector(7 downto 0);
    signal IMC19_8862 : std_logic_vector(7 downto 0);
    signal IMC1_8718 : std_logic_vector(7 downto 0);
    signal IMC20_8870 : std_logic_vector(7 downto 0);
    signal IMC21_8878 : std_logic_vector(7 downto 0);
    signal IMC22_8886 : std_logic_vector(7 downto 0);
    signal IMC23_8894 : std_logic_vector(7 downto 0);
    signal IMC24_8902 : std_logic_vector(7 downto 0);
    signal IMC25_8910 : std_logic_vector(7 downto 0);
    signal IMC26_8918 : std_logic_vector(7 downto 0);
    signal IMC27_8926 : std_logic_vector(7 downto 0);
    signal IMC28_8934 : std_logic_vector(7 downto 0);
    signal IMC29_8942 : std_logic_vector(7 downto 0);
    signal IMC2_8726 : std_logic_vector(7 downto 0);
    signal IMC30_8950 : std_logic_vector(7 downto 0);
    signal IMC31_8958 : std_logic_vector(7 downto 0);
    signal IMC3_8734 : std_logic_vector(7 downto 0);
    signal IMC4_8742 : std_logic_vector(7 downto 0);
    signal IMC5_8750 : std_logic_vector(7 downto 0);
    signal IMC6_8758 : std_logic_vector(7 downto 0);
    signal IMC7_8766 : std_logic_vector(7 downto 0);
    signal IMC8_8774 : std_logic_vector(7 downto 0);
    signal IMC9_8782 : std_logic_vector(7 downto 0);
    signal IMD0_8966 : std_logic_vector(7 downto 0);
    signal IMD10_9046 : std_logic_vector(7 downto 0);
    signal IMD11_9054 : std_logic_vector(7 downto 0);
    signal IMD12_9062 : std_logic_vector(7 downto 0);
    signal IMD13_9070 : std_logic_vector(7 downto 0);
    signal IMD14_9078 : std_logic_vector(7 downto 0);
    signal IMD15_9086 : std_logic_vector(7 downto 0);
    signal IMD1_8974 : std_logic_vector(7 downto 0);
    signal IMD2_8982 : std_logic_vector(7 downto 0);
    signal IMD3_8990 : std_logic_vector(7 downto 0);
    signal IMD4_8998 : std_logic_vector(7 downto 0);
    signal IMD5_9006 : std_logic_vector(7 downto 0);
    signal IMD6_9014 : std_logic_vector(7 downto 0);
    signal IMD7_9022 : std_logic_vector(7 downto 0);
    signal IMD8_9030 : std_logic_vector(7 downto 0);
    signal IMD9_9038 : std_logic_vector(7 downto 0);
    signal IME0_9094 : std_logic_vector(7 downto 0);
    signal IME1_9102 : std_logic_vector(7 downto 0);
    signal IME2_9110 : std_logic_vector(7 downto 0);
    signal IME3_9118 : std_logic_vector(7 downto 0);
    signal IME4_9126 : std_logic_vector(7 downto 0);
    signal IME5_9134 : std_logic_vector(7 downto 0);
    signal IME6_9142 : std_logic_vector(7 downto 0);
    signal IME7_9150 : std_logic_vector(7 downto 0);
    signal IMF0_9158 : std_logic_vector(7 downto 0);
    signal IMF1_9166 : std_logic_vector(7 downto 0);
    signal IMF2_9174 : std_logic_vector(7 downto 0);
    signal IMF3_9182 : std_logic_vector(7 downto 0);
    signal IMG0_9190 : std_logic_vector(7 downto 0);
    signal IMG1_9198 : std_logic_vector(7 downto 0);
    signal konst_6913_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6923_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6933_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6943_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6953_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6963_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6973_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6983_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6993_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7003_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7013_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7023_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7033_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7043_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7053_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7063_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7073_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7083_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7093_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7103_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7113_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7123_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7133_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7143_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7153_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7163_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7173_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7183_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7193_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7203_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7213_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7223_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7233_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7243_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7253_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7263_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7273_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7283_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7293_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7303_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7313_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7323_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7333_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7343_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7353_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7363_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7373_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7383_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7393_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7403_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7413_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7423_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7433_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7443_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7453_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7463_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7473_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7483_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7493_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7503_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7513_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7523_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7533_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7543_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7553_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7563_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7573_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7583_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7593_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7603_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7613_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7623_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7633_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7643_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7653_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7663_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7673_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7683_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7693_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7703_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7713_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7723_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7733_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7743_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7753_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7763_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7773_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7783_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7793_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7803_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7813_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7823_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7833_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7843_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7853_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7863_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7873_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7883_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7893_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7903_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7913_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7923_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7933_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7943_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7953_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7963_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7973_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7983_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7993_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8003_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8013_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8023_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8033_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8043_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8053_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8063_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8073_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8083_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8093_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8103_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8113_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8123_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8133_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8143_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8153_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8163_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8173_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8183_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8193_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8201_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8209_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8217_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8225_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8233_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8241_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8249_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8257_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8265_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8273_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8281_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8289_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8297_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8305_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8313_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8321_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8329_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8337_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8345_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8353_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8361_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8369_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8377_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8385_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8393_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8401_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8409_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8417_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8425_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8433_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8441_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8449_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8457_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8465_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8473_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8481_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8489_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8497_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8505_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8513_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8521_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8529_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8537_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8545_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8553_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8561_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8569_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8577_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8585_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8593_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8601_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8609_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8617_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8625_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8633_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8641_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8649_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8657_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8665_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8673_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8681_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8689_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8697_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8705_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8713_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8721_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8729_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8737_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8745_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8753_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8761_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8769_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8777_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8785_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8793_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8801_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8809_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8817_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8825_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8833_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8841_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8849_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8857_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8865_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8873_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8881_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8889_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8897_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8905_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8913_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8921_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8929_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8937_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8945_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8953_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8961_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8969_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8977_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8985_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8993_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9001_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9009_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9017_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9025_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9033_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9041_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9049_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9057_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9065_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9073_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9081_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9089_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9097_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9105_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9113_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9121_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9129_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9137_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9145_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9153_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9161_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9169_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9177_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9185_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9193_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9201_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_6916_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_6918_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_6926_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_6928_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_6936_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_6938_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_6946_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_6948_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_6956_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_6958_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_6966_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_6968_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_6976_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_6978_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_6986_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_6988_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_6996_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_6998_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7006_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7008_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7016_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7018_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7026_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7028_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7036_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7038_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7046_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7048_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7056_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7058_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7066_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7068_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7076_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7078_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7086_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7088_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7096_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7098_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7106_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7108_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7116_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7118_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7126_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7128_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7136_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7138_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7146_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7148_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7156_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7158_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7166_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7168_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7176_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7178_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7186_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7188_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7196_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7198_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7206_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7208_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7216_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7218_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7226_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7228_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7236_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7238_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7246_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7248_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7256_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7258_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7266_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7268_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7276_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7278_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7286_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7288_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7296_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7298_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7306_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7308_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7316_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7318_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7326_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7328_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7336_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7338_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7346_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7348_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7356_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7358_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7366_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7368_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7376_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7378_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7386_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7388_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7396_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7398_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7406_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7408_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7416_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7418_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7426_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7428_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7436_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7438_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7446_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7448_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7456_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7458_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7466_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7468_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7476_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7478_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7486_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7488_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7496_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7498_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7506_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7508_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7516_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7518_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7526_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7528_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7536_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7538_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7546_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7548_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7556_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7558_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7566_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7568_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7576_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7578_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7586_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7588_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7596_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7598_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7606_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7608_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7616_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7618_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7626_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7628_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7636_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7638_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7646_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7648_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7656_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7658_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7666_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7668_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7676_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7678_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7686_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7688_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7696_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7698_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7706_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7708_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7716_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7718_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7726_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7728_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7736_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7738_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7746_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7748_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7756_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7758_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7766_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7768_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7776_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7778_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7786_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7788_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7796_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7798_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7806_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7808_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7816_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7818_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7826_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7828_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7836_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7838_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7846_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7848_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7856_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7858_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7866_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7868_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7876_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7878_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7886_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7888_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7896_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7898_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7906_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7908_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7916_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7918_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7926_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7928_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7936_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7938_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7946_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7948_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7956_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7958_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7966_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7968_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7976_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7978_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7986_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7988_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7996_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7998_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_8006_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_8008_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_8016_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_8018_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_8026_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_8028_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_8036_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_8038_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_8046_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_8048_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_8056_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_8058_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_8066_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_8068_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_8076_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_8078_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_8086_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_8088_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_8096_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_8098_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_8106_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_8108_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_8116_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_8118_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_8126_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_8128_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_8136_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_8138_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_8146_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_8148_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_8156_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_8158_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_8166_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_8168_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_8176_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_8178_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_8186_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_8188_wire_constant : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    konst_6913_wire_constant <= "00000000";
    konst_6923_wire_constant <= "00000000";
    konst_6933_wire_constant <= "00000000";
    konst_6943_wire_constant <= "00000000";
    konst_6953_wire_constant <= "00000000";
    konst_6963_wire_constant <= "00000000";
    konst_6973_wire_constant <= "00000000";
    konst_6983_wire_constant <= "00000000";
    konst_6993_wire_constant <= "00000000";
    konst_7003_wire_constant <= "00000000";
    konst_7013_wire_constant <= "00000000";
    konst_7023_wire_constant <= "00000000";
    konst_7033_wire_constant <= "00000000";
    konst_7043_wire_constant <= "00000000";
    konst_7053_wire_constant <= "00000000";
    konst_7063_wire_constant <= "00000000";
    konst_7073_wire_constant <= "00000000";
    konst_7083_wire_constant <= "00000000";
    konst_7093_wire_constant <= "00000000";
    konst_7103_wire_constant <= "00000000";
    konst_7113_wire_constant <= "00000000";
    konst_7123_wire_constant <= "00000000";
    konst_7133_wire_constant <= "00000000";
    konst_7143_wire_constant <= "00000000";
    konst_7153_wire_constant <= "00000000";
    konst_7163_wire_constant <= "00000000";
    konst_7173_wire_constant <= "00000000";
    konst_7183_wire_constant <= "00000000";
    konst_7193_wire_constant <= "00000000";
    konst_7203_wire_constant <= "00000000";
    konst_7213_wire_constant <= "00000000";
    konst_7223_wire_constant <= "00000000";
    konst_7233_wire_constant <= "00000000";
    konst_7243_wire_constant <= "00000000";
    konst_7253_wire_constant <= "00000000";
    konst_7263_wire_constant <= "00000000";
    konst_7273_wire_constant <= "00000000";
    konst_7283_wire_constant <= "00000000";
    konst_7293_wire_constant <= "00000000";
    konst_7303_wire_constant <= "00000000";
    konst_7313_wire_constant <= "00000000";
    konst_7323_wire_constant <= "00000000";
    konst_7333_wire_constant <= "00000000";
    konst_7343_wire_constant <= "00000000";
    konst_7353_wire_constant <= "00000000";
    konst_7363_wire_constant <= "00000000";
    konst_7373_wire_constant <= "00000000";
    konst_7383_wire_constant <= "00000000";
    konst_7393_wire_constant <= "00000000";
    konst_7403_wire_constant <= "00000000";
    konst_7413_wire_constant <= "00000000";
    konst_7423_wire_constant <= "00000000";
    konst_7433_wire_constant <= "00000000";
    konst_7443_wire_constant <= "00000000";
    konst_7453_wire_constant <= "00000000";
    konst_7463_wire_constant <= "00000000";
    konst_7473_wire_constant <= "00000000";
    konst_7483_wire_constant <= "00000000";
    konst_7493_wire_constant <= "00000000";
    konst_7503_wire_constant <= "00000000";
    konst_7513_wire_constant <= "00000000";
    konst_7523_wire_constant <= "00000000";
    konst_7533_wire_constant <= "00000000";
    konst_7543_wire_constant <= "00000000";
    konst_7553_wire_constant <= "00000000";
    konst_7563_wire_constant <= "00000000";
    konst_7573_wire_constant <= "00000000";
    konst_7583_wire_constant <= "00000000";
    konst_7593_wire_constant <= "00000000";
    konst_7603_wire_constant <= "00000000";
    konst_7613_wire_constant <= "00000000";
    konst_7623_wire_constant <= "00000000";
    konst_7633_wire_constant <= "00000000";
    konst_7643_wire_constant <= "00000000";
    konst_7653_wire_constant <= "00000000";
    konst_7663_wire_constant <= "00000000";
    konst_7673_wire_constant <= "00000000";
    konst_7683_wire_constant <= "00000000";
    konst_7693_wire_constant <= "00000000";
    konst_7703_wire_constant <= "00000000";
    konst_7713_wire_constant <= "00000000";
    konst_7723_wire_constant <= "00000000";
    konst_7733_wire_constant <= "00000000";
    konst_7743_wire_constant <= "00000000";
    konst_7753_wire_constant <= "00000000";
    konst_7763_wire_constant <= "00000000";
    konst_7773_wire_constant <= "00000000";
    konst_7783_wire_constant <= "00000000";
    konst_7793_wire_constant <= "00000000";
    konst_7803_wire_constant <= "00000000";
    konst_7813_wire_constant <= "00000000";
    konst_7823_wire_constant <= "00000000";
    konst_7833_wire_constant <= "00000000";
    konst_7843_wire_constant <= "00000000";
    konst_7853_wire_constant <= "00000000";
    konst_7863_wire_constant <= "00000000";
    konst_7873_wire_constant <= "00000000";
    konst_7883_wire_constant <= "00000000";
    konst_7893_wire_constant <= "00000000";
    konst_7903_wire_constant <= "00000000";
    konst_7913_wire_constant <= "00000000";
    konst_7923_wire_constant <= "00000000";
    konst_7933_wire_constant <= "00000000";
    konst_7943_wire_constant <= "00000000";
    konst_7953_wire_constant <= "00000000";
    konst_7963_wire_constant <= "00000000";
    konst_7973_wire_constant <= "00000000";
    konst_7983_wire_constant <= "00000000";
    konst_7993_wire_constant <= "00000000";
    konst_8003_wire_constant <= "00000000";
    konst_8013_wire_constant <= "00000000";
    konst_8023_wire_constant <= "00000000";
    konst_8033_wire_constant <= "00000000";
    konst_8043_wire_constant <= "00000000";
    konst_8053_wire_constant <= "00000000";
    konst_8063_wire_constant <= "00000000";
    konst_8073_wire_constant <= "00000000";
    konst_8083_wire_constant <= "00000000";
    konst_8093_wire_constant <= "00000000";
    konst_8103_wire_constant <= "00000000";
    konst_8113_wire_constant <= "00000000";
    konst_8123_wire_constant <= "00000000";
    konst_8133_wire_constant <= "00000000";
    konst_8143_wire_constant <= "00000000";
    konst_8153_wire_constant <= "00000000";
    konst_8163_wire_constant <= "00000000";
    konst_8173_wire_constant <= "00000000";
    konst_8183_wire_constant <= "00000000";
    konst_8193_wire_constant <= "00000001";
    konst_8201_wire_constant <= "00000001";
    konst_8209_wire_constant <= "00000001";
    konst_8217_wire_constant <= "00000001";
    konst_8225_wire_constant <= "00000001";
    konst_8233_wire_constant <= "00000001";
    konst_8241_wire_constant <= "00000001";
    konst_8249_wire_constant <= "00000001";
    konst_8257_wire_constant <= "00000001";
    konst_8265_wire_constant <= "00000001";
    konst_8273_wire_constant <= "00000001";
    konst_8281_wire_constant <= "00000001";
    konst_8289_wire_constant <= "00000001";
    konst_8297_wire_constant <= "00000001";
    konst_8305_wire_constant <= "00000001";
    konst_8313_wire_constant <= "00000001";
    konst_8321_wire_constant <= "00000001";
    konst_8329_wire_constant <= "00000001";
    konst_8337_wire_constant <= "00000001";
    konst_8345_wire_constant <= "00000001";
    konst_8353_wire_constant <= "00000001";
    konst_8361_wire_constant <= "00000001";
    konst_8369_wire_constant <= "00000001";
    konst_8377_wire_constant <= "00000001";
    konst_8385_wire_constant <= "00000001";
    konst_8393_wire_constant <= "00000001";
    konst_8401_wire_constant <= "00000001";
    konst_8409_wire_constant <= "00000001";
    konst_8417_wire_constant <= "00000001";
    konst_8425_wire_constant <= "00000001";
    konst_8433_wire_constant <= "00000001";
    konst_8441_wire_constant <= "00000001";
    konst_8449_wire_constant <= "00000001";
    konst_8457_wire_constant <= "00000001";
    konst_8465_wire_constant <= "00000001";
    konst_8473_wire_constant <= "00000001";
    konst_8481_wire_constant <= "00000001";
    konst_8489_wire_constant <= "00000001";
    konst_8497_wire_constant <= "00000001";
    konst_8505_wire_constant <= "00000001";
    konst_8513_wire_constant <= "00000001";
    konst_8521_wire_constant <= "00000001";
    konst_8529_wire_constant <= "00000001";
    konst_8537_wire_constant <= "00000001";
    konst_8545_wire_constant <= "00000001";
    konst_8553_wire_constant <= "00000001";
    konst_8561_wire_constant <= "00000001";
    konst_8569_wire_constant <= "00000001";
    konst_8577_wire_constant <= "00000001";
    konst_8585_wire_constant <= "00000001";
    konst_8593_wire_constant <= "00000001";
    konst_8601_wire_constant <= "00000001";
    konst_8609_wire_constant <= "00000001";
    konst_8617_wire_constant <= "00000001";
    konst_8625_wire_constant <= "00000001";
    konst_8633_wire_constant <= "00000001";
    konst_8641_wire_constant <= "00000001";
    konst_8649_wire_constant <= "00000001";
    konst_8657_wire_constant <= "00000001";
    konst_8665_wire_constant <= "00000001";
    konst_8673_wire_constant <= "00000001";
    konst_8681_wire_constant <= "00000001";
    konst_8689_wire_constant <= "00000001";
    konst_8697_wire_constant <= "00000001";
    konst_8705_wire_constant <= "00000010";
    konst_8713_wire_constant <= "00000010";
    konst_8721_wire_constant <= "00000010";
    konst_8729_wire_constant <= "00000010";
    konst_8737_wire_constant <= "00000010";
    konst_8745_wire_constant <= "00000010";
    konst_8753_wire_constant <= "00000010";
    konst_8761_wire_constant <= "00000010";
    konst_8769_wire_constant <= "00000010";
    konst_8777_wire_constant <= "00000010";
    konst_8785_wire_constant <= "00000010";
    konst_8793_wire_constant <= "00000010";
    konst_8801_wire_constant <= "00000010";
    konst_8809_wire_constant <= "00000010";
    konst_8817_wire_constant <= "00000010";
    konst_8825_wire_constant <= "00000010";
    konst_8833_wire_constant <= "00000010";
    konst_8841_wire_constant <= "00000010";
    konst_8849_wire_constant <= "00000010";
    konst_8857_wire_constant <= "00000010";
    konst_8865_wire_constant <= "00000010";
    konst_8873_wire_constant <= "00000010";
    konst_8881_wire_constant <= "00000010";
    konst_8889_wire_constant <= "00000010";
    konst_8897_wire_constant <= "00000010";
    konst_8905_wire_constant <= "00000010";
    konst_8913_wire_constant <= "00000010";
    konst_8921_wire_constant <= "00000010";
    konst_8929_wire_constant <= "00000010";
    konst_8937_wire_constant <= "00000010";
    konst_8945_wire_constant <= "00000010";
    konst_8953_wire_constant <= "00000010";
    konst_8961_wire_constant <= "00000011";
    konst_8969_wire_constant <= "00000011";
    konst_8977_wire_constant <= "00000011";
    konst_8985_wire_constant <= "00000011";
    konst_8993_wire_constant <= "00000011";
    konst_9001_wire_constant <= "00000011";
    konst_9009_wire_constant <= "00000011";
    konst_9017_wire_constant <= "00000011";
    konst_9025_wire_constant <= "00000011";
    konst_9033_wire_constant <= "00000011";
    konst_9041_wire_constant <= "00000011";
    konst_9049_wire_constant <= "00000011";
    konst_9057_wire_constant <= "00000011";
    konst_9065_wire_constant <= "00000011";
    konst_9073_wire_constant <= "00000011";
    konst_9081_wire_constant <= "00000011";
    konst_9089_wire_constant <= "00000100";
    konst_9097_wire_constant <= "00000100";
    konst_9105_wire_constant <= "00000100";
    konst_9113_wire_constant <= "00000100";
    konst_9121_wire_constant <= "00000100";
    konst_9129_wire_constant <= "00000100";
    konst_9137_wire_constant <= "00000100";
    konst_9145_wire_constant <= "00000100";
    konst_9153_wire_constant <= "00000101";
    konst_9161_wire_constant <= "00000101";
    konst_9169_wire_constant <= "00000101";
    konst_9177_wire_constant <= "00000101";
    konst_9185_wire_constant <= "00000110";
    konst_9193_wire_constant <= "00000110";
    konst_9201_wire_constant <= "00000111";
    type_cast_6916_wire_constant <= "00001001";
    type_cast_6918_wire_constant <= "01010010";
    type_cast_6926_wire_constant <= "11010101";
    type_cast_6928_wire_constant <= "01101010";
    type_cast_6936_wire_constant <= "00110110";
    type_cast_6938_wire_constant <= "00110000";
    type_cast_6946_wire_constant <= "00111000";
    type_cast_6948_wire_constant <= "10100101";
    type_cast_6956_wire_constant <= "01000000";
    type_cast_6958_wire_constant <= "10111111";
    type_cast_6966_wire_constant <= "10011110";
    type_cast_6968_wire_constant <= "10100011";
    type_cast_6976_wire_constant <= "11110011";
    type_cast_6978_wire_constant <= "10000001";
    type_cast_6986_wire_constant <= "11111011";
    type_cast_6988_wire_constant <= "11010111";
    type_cast_6996_wire_constant <= "11100011";
    type_cast_6998_wire_constant <= "01111100";
    type_cast_7006_wire_constant <= "10000010";
    type_cast_7008_wire_constant <= "00111001";
    type_cast_7016_wire_constant <= "00101111";
    type_cast_7018_wire_constant <= "10011011";
    type_cast_7026_wire_constant <= "10000111";
    type_cast_7028_wire_constant <= "11111111";
    type_cast_7036_wire_constant <= "10001110";
    type_cast_7038_wire_constant <= "00110100";
    type_cast_7046_wire_constant <= "01000100";
    type_cast_7048_wire_constant <= "01000011";
    type_cast_7056_wire_constant <= "11011110";
    type_cast_7058_wire_constant <= "11000100";
    type_cast_7066_wire_constant <= "11001011";
    type_cast_7068_wire_constant <= "11101001";
    type_cast_7076_wire_constant <= "01111011";
    type_cast_7078_wire_constant <= "01010100";
    type_cast_7086_wire_constant <= "00110010";
    type_cast_7088_wire_constant <= "10010100";
    type_cast_7096_wire_constant <= "11000010";
    type_cast_7098_wire_constant <= "10100110";
    type_cast_7106_wire_constant <= "00111101";
    type_cast_7108_wire_constant <= "00100011";
    type_cast_7116_wire_constant <= "01001100";
    type_cast_7118_wire_constant <= "11101110";
    type_cast_7126_wire_constant <= "00001011";
    type_cast_7128_wire_constant <= "10010101";
    type_cast_7136_wire_constant <= "11111010";
    type_cast_7138_wire_constant <= "01000010";
    type_cast_7146_wire_constant <= "01001110";
    type_cast_7148_wire_constant <= "11000011";
    type_cast_7156_wire_constant <= "00101110";
    type_cast_7158_wire_constant <= "00001000";
    type_cast_7166_wire_constant <= "01100110";
    type_cast_7168_wire_constant <= "10100001";
    type_cast_7176_wire_constant <= "11011001";
    type_cast_7178_wire_constant <= "00101000";
    type_cast_7186_wire_constant <= "10110010";
    type_cast_7188_wire_constant <= "00100100";
    type_cast_7196_wire_constant <= "01011011";
    type_cast_7198_wire_constant <= "01110110";
    type_cast_7206_wire_constant <= "01001001";
    type_cast_7208_wire_constant <= "10100010";
    type_cast_7216_wire_constant <= "10001011";
    type_cast_7218_wire_constant <= "01101101";
    type_cast_7226_wire_constant <= "00100101";
    type_cast_7228_wire_constant <= "11010001";
    type_cast_7236_wire_constant <= "11111000";
    type_cast_7238_wire_constant <= "01110010";
    type_cast_7246_wire_constant <= "01100100";
    type_cast_7248_wire_constant <= "11110110";
    type_cast_7256_wire_constant <= "01101000";
    type_cast_7258_wire_constant <= "10000110";
    type_cast_7266_wire_constant <= "00010110";
    type_cast_7268_wire_constant <= "10011000";
    type_cast_7276_wire_constant <= "10100100";
    type_cast_7278_wire_constant <= "11010100";
    type_cast_7286_wire_constant <= "11001100";
    type_cast_7288_wire_constant <= "01011100";
    type_cast_7296_wire_constant <= "01100101";
    type_cast_7298_wire_constant <= "01011101";
    type_cast_7306_wire_constant <= "10010010";
    type_cast_7308_wire_constant <= "10110110";
    type_cast_7316_wire_constant <= "01110000";
    type_cast_7318_wire_constant <= "01101100";
    type_cast_7326_wire_constant <= "01010000";
    type_cast_7328_wire_constant <= "01001000";
    type_cast_7336_wire_constant <= "11101101";
    type_cast_7338_wire_constant <= "11111101";
    type_cast_7346_wire_constant <= "11011010";
    type_cast_7348_wire_constant <= "10111001";
    type_cast_7356_wire_constant <= "00010101";
    type_cast_7358_wire_constant <= "01011110";
    type_cast_7366_wire_constant <= "01010111";
    type_cast_7368_wire_constant <= "01000110";
    type_cast_7376_wire_constant <= "10001101";
    type_cast_7378_wire_constant <= "10100111";
    type_cast_7386_wire_constant <= "10000100";
    type_cast_7388_wire_constant <= "10011101";
    type_cast_7396_wire_constant <= "11011000";
    type_cast_7398_wire_constant <= "10010000";
    type_cast_7406_wire_constant <= "00000000";
    type_cast_7408_wire_constant <= "10101011";
    type_cast_7416_wire_constant <= "10111100";
    type_cast_7418_wire_constant <= "10001100";
    type_cast_7426_wire_constant <= "00001010";
    type_cast_7428_wire_constant <= "11010011";
    type_cast_7436_wire_constant <= "11100100";
    type_cast_7438_wire_constant <= "11110111";
    type_cast_7446_wire_constant <= "00000101";
    type_cast_7448_wire_constant <= "01011000";
    type_cast_7456_wire_constant <= "10110011";
    type_cast_7458_wire_constant <= "10111000";
    type_cast_7466_wire_constant <= "00000110";
    type_cast_7468_wire_constant <= "01000101";
    type_cast_7476_wire_constant <= "00101100";
    type_cast_7478_wire_constant <= "11010000";
    type_cast_7486_wire_constant <= "10001111";
    type_cast_7488_wire_constant <= "00011110";
    type_cast_7496_wire_constant <= "00111111";
    type_cast_7498_wire_constant <= "11001010";
    type_cast_7506_wire_constant <= "00000010";
    type_cast_7508_wire_constant <= "00001111";
    type_cast_7516_wire_constant <= "10101111";
    type_cast_7518_wire_constant <= "11000001";
    type_cast_7526_wire_constant <= "00000011";
    type_cast_7528_wire_constant <= "10111101";
    type_cast_7536_wire_constant <= "00010011";
    type_cast_7538_wire_constant <= "00000001";
    type_cast_7546_wire_constant <= "01101011";
    type_cast_7548_wire_constant <= "10001010";
    type_cast_7556_wire_constant <= "10010001";
    type_cast_7558_wire_constant <= "00111010";
    type_cast_7566_wire_constant <= "01000001";
    type_cast_7568_wire_constant <= "00010001";
    type_cast_7576_wire_constant <= "01100111";
    type_cast_7578_wire_constant <= "01001111";
    type_cast_7586_wire_constant <= "11101010";
    type_cast_7588_wire_constant <= "11011100";
    type_cast_7596_wire_constant <= "11110010";
    type_cast_7598_wire_constant <= "10010111";
    type_cast_7606_wire_constant <= "11001110";
    type_cast_7608_wire_constant <= "11001111";
    type_cast_7616_wire_constant <= "10110100";
    type_cast_7618_wire_constant <= "11110000";
    type_cast_7626_wire_constant <= "01110011";
    type_cast_7628_wire_constant <= "11100110";
    type_cast_7636_wire_constant <= "10101100";
    type_cast_7638_wire_constant <= "10010110";
    type_cast_7646_wire_constant <= "00100010";
    type_cast_7648_wire_constant <= "01110100";
    type_cast_7656_wire_constant <= "10101101";
    type_cast_7658_wire_constant <= "11100111";
    type_cast_7666_wire_constant <= "10000101";
    type_cast_7668_wire_constant <= "00110101";
    type_cast_7676_wire_constant <= "11111001";
    type_cast_7678_wire_constant <= "11100010";
    type_cast_7686_wire_constant <= "11101000";
    type_cast_7688_wire_constant <= "00110111";
    type_cast_7696_wire_constant <= "01110101";
    type_cast_7698_wire_constant <= "00011100";
    type_cast_7706_wire_constant <= "01101110";
    type_cast_7708_wire_constant <= "11011111";
    type_cast_7716_wire_constant <= "11110001";
    type_cast_7718_wire_constant <= "01000111";
    type_cast_7726_wire_constant <= "01110001";
    type_cast_7728_wire_constant <= "00011010";
    type_cast_7736_wire_constant <= "00101001";
    type_cast_7738_wire_constant <= "00011101";
    type_cast_7746_wire_constant <= "10001001";
    type_cast_7748_wire_constant <= "11000101";
    type_cast_7756_wire_constant <= "10110111";
    type_cast_7758_wire_constant <= "01101111";
    type_cast_7766_wire_constant <= "00001110";
    type_cast_7768_wire_constant <= "01100010";
    type_cast_7776_wire_constant <= "00011000";
    type_cast_7778_wire_constant <= "10101010";
    type_cast_7786_wire_constant <= "00011011";
    type_cast_7788_wire_constant <= "10111110";
    type_cast_7796_wire_constant <= "01010110";
    type_cast_7798_wire_constant <= "11111100";
    type_cast_7806_wire_constant <= "01001011";
    type_cast_7808_wire_constant <= "00111110";
    type_cast_7816_wire_constant <= "11010010";
    type_cast_7818_wire_constant <= "11000110";
    type_cast_7826_wire_constant <= "00100000";
    type_cast_7828_wire_constant <= "01111001";
    type_cast_7836_wire_constant <= "11011011";
    type_cast_7838_wire_constant <= "10011010";
    type_cast_7846_wire_constant <= "11111110";
    type_cast_7848_wire_constant <= "11000000";
    type_cast_7856_wire_constant <= "11001101";
    type_cast_7858_wire_constant <= "01111000";
    type_cast_7866_wire_constant <= "11110100";
    type_cast_7868_wire_constant <= "01011010";
    type_cast_7876_wire_constant <= "11011101";
    type_cast_7878_wire_constant <= "00011111";
    type_cast_7886_wire_constant <= "00110011";
    type_cast_7888_wire_constant <= "10101000";
    type_cast_7896_wire_constant <= "00000111";
    type_cast_7898_wire_constant <= "10001000";
    type_cast_7906_wire_constant <= "00110001";
    type_cast_7908_wire_constant <= "11000111";
    type_cast_7916_wire_constant <= "00010010";
    type_cast_7918_wire_constant <= "10110001";
    type_cast_7926_wire_constant <= "01011001";
    type_cast_7928_wire_constant <= "00010000";
    type_cast_7936_wire_constant <= "10000000";
    type_cast_7938_wire_constant <= "00100111";
    type_cast_7946_wire_constant <= "01011111";
    type_cast_7948_wire_constant <= "11101100";
    type_cast_7956_wire_constant <= "01010001";
    type_cast_7958_wire_constant <= "01100000";
    type_cast_7966_wire_constant <= "10101001";
    type_cast_7968_wire_constant <= "01111111";
    type_cast_7976_wire_constant <= "10110101";
    type_cast_7978_wire_constant <= "00011001";
    type_cast_7986_wire_constant <= "00001101";
    type_cast_7988_wire_constant <= "01001010";
    type_cast_7996_wire_constant <= "11100101";
    type_cast_7998_wire_constant <= "00101101";
    type_cast_8006_wire_constant <= "10011111";
    type_cast_8008_wire_constant <= "01111010";
    type_cast_8016_wire_constant <= "11001001";
    type_cast_8018_wire_constant <= "10010011";
    type_cast_8026_wire_constant <= "11101111";
    type_cast_8028_wire_constant <= "10011100";
    type_cast_8036_wire_constant <= "11100000";
    type_cast_8038_wire_constant <= "10100000";
    type_cast_8046_wire_constant <= "01001101";
    type_cast_8048_wire_constant <= "00111011";
    type_cast_8056_wire_constant <= "00101010";
    type_cast_8058_wire_constant <= "10101110";
    type_cast_8066_wire_constant <= "10110000";
    type_cast_8068_wire_constant <= "11110101";
    type_cast_8076_wire_constant <= "11101011";
    type_cast_8078_wire_constant <= "11001000";
    type_cast_8086_wire_constant <= "00111100";
    type_cast_8088_wire_constant <= "10111011";
    type_cast_8096_wire_constant <= "01010011";
    type_cast_8098_wire_constant <= "10000011";
    type_cast_8106_wire_constant <= "01100001";
    type_cast_8108_wire_constant <= "10011001";
    type_cast_8116_wire_constant <= "00101011";
    type_cast_8118_wire_constant <= "00010111";
    type_cast_8126_wire_constant <= "01111110";
    type_cast_8128_wire_constant <= "00000100";
    type_cast_8136_wire_constant <= "01110111";
    type_cast_8138_wire_constant <= "10111010";
    type_cast_8146_wire_constant <= "00100110";
    type_cast_8148_wire_constant <= "11010110";
    type_cast_8156_wire_constant <= "01101001";
    type_cast_8158_wire_constant <= "11100001";
    type_cast_8166_wire_constant <= "01100011";
    type_cast_8168_wire_constant <= "00010100";
    type_cast_8176_wire_constant <= "00100001";
    type_cast_8178_wire_constant <= "01010101";
    type_cast_8186_wire_constant <= "01111101";
    type_cast_8188_wire_constant <= "00001100";
    -- logger for split-operator MUX_6919_inst flow-through 
    process(IMA0_6920) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_6919_inst:flowthrough inputs: " & " BITSEL_u8_u1_6914_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6914_wire) & " type_cast_6916_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_6916_wire_constant) & " type_cast_6918_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_6918_wire_constant) & " outputs:" & " IMA0_6920= "  & Convert_SLV_To_Hex_String(IMA0_6920));
      --
    end process; 
    -- flow-through select operator MUX_6919_inst
    IMA0_6920 <= type_cast_6916_wire_constant when (BITSEL_u8_u1_6914_wire(0) /=  '0') else type_cast_6918_wire_constant;
    -- logger for split-operator MUX_6929_inst flow-through 
    process(IMA1_6930) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_6929_inst:flowthrough inputs: " & " BITSEL_u8_u1_6924_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6924_wire) & " type_cast_6926_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_6926_wire_constant) & " type_cast_6928_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_6928_wire_constant) & " outputs:" & " IMA1_6930= "  & Convert_SLV_To_Hex_String(IMA1_6930));
      --
    end process; 
    -- flow-through select operator MUX_6929_inst
    IMA1_6930 <= type_cast_6926_wire_constant when (BITSEL_u8_u1_6924_wire(0) /=  '0') else type_cast_6928_wire_constant;
    -- logger for split-operator MUX_6939_inst flow-through 
    process(IMA2_6940) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_6939_inst:flowthrough inputs: " & " BITSEL_u8_u1_6934_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6934_wire) & " type_cast_6936_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_6936_wire_constant) & " type_cast_6938_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_6938_wire_constant) & " outputs:" & " IMA2_6940= "  & Convert_SLV_To_Hex_String(IMA2_6940));
      --
    end process; 
    -- flow-through select operator MUX_6939_inst
    IMA2_6940 <= type_cast_6936_wire_constant when (BITSEL_u8_u1_6934_wire(0) /=  '0') else type_cast_6938_wire_constant;
    -- logger for split-operator MUX_6949_inst flow-through 
    process(IMA3_6950) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_6949_inst:flowthrough inputs: " & " BITSEL_u8_u1_6944_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6944_wire) & " type_cast_6946_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_6946_wire_constant) & " type_cast_6948_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_6948_wire_constant) & " outputs:" & " IMA3_6950= "  & Convert_SLV_To_Hex_String(IMA3_6950));
      --
    end process; 
    -- flow-through select operator MUX_6949_inst
    IMA3_6950 <= type_cast_6946_wire_constant when (BITSEL_u8_u1_6944_wire(0) /=  '0') else type_cast_6948_wire_constant;
    -- logger for split-operator MUX_6959_inst flow-through 
    process(IMA4_6960) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_6959_inst:flowthrough inputs: " & " BITSEL_u8_u1_6954_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6954_wire) & " type_cast_6956_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_6956_wire_constant) & " type_cast_6958_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_6958_wire_constant) & " outputs:" & " IMA4_6960= "  & Convert_SLV_To_Hex_String(IMA4_6960));
      --
    end process; 
    -- flow-through select operator MUX_6959_inst
    IMA4_6960 <= type_cast_6956_wire_constant when (BITSEL_u8_u1_6954_wire(0) /=  '0') else type_cast_6958_wire_constant;
    -- logger for split-operator MUX_6969_inst flow-through 
    process(IMA5_6970) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_6969_inst:flowthrough inputs: " & " BITSEL_u8_u1_6964_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6964_wire) & " type_cast_6966_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_6966_wire_constant) & " type_cast_6968_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_6968_wire_constant) & " outputs:" & " IMA5_6970= "  & Convert_SLV_To_Hex_String(IMA5_6970));
      --
    end process; 
    -- flow-through select operator MUX_6969_inst
    IMA5_6970 <= type_cast_6966_wire_constant when (BITSEL_u8_u1_6964_wire(0) /=  '0') else type_cast_6968_wire_constant;
    -- logger for split-operator MUX_6979_inst flow-through 
    process(IMA6_6980) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_6979_inst:flowthrough inputs: " & " BITSEL_u8_u1_6974_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6974_wire) & " type_cast_6976_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_6976_wire_constant) & " type_cast_6978_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_6978_wire_constant) & " outputs:" & " IMA6_6980= "  & Convert_SLV_To_Hex_String(IMA6_6980));
      --
    end process; 
    -- flow-through select operator MUX_6979_inst
    IMA6_6980 <= type_cast_6976_wire_constant when (BITSEL_u8_u1_6974_wire(0) /=  '0') else type_cast_6978_wire_constant;
    -- logger for split-operator MUX_6989_inst flow-through 
    process(IMA7_6990) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_6989_inst:flowthrough inputs: " & " BITSEL_u8_u1_6984_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6984_wire) & " type_cast_6986_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_6986_wire_constant) & " type_cast_6988_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_6988_wire_constant) & " outputs:" & " IMA7_6990= "  & Convert_SLV_To_Hex_String(IMA7_6990));
      --
    end process; 
    -- flow-through select operator MUX_6989_inst
    IMA7_6990 <= type_cast_6986_wire_constant when (BITSEL_u8_u1_6984_wire(0) /=  '0') else type_cast_6988_wire_constant;
    -- logger for split-operator MUX_6999_inst flow-through 
    process(IMA8_7000) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_6999_inst:flowthrough inputs: " & " BITSEL_u8_u1_6994_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_6994_wire) & " type_cast_6996_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_6996_wire_constant) & " type_cast_6998_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_6998_wire_constant) & " outputs:" & " IMA8_7000= "  & Convert_SLV_To_Hex_String(IMA8_7000));
      --
    end process; 
    -- flow-through select operator MUX_6999_inst
    IMA8_7000 <= type_cast_6996_wire_constant when (BITSEL_u8_u1_6994_wire(0) /=  '0') else type_cast_6998_wire_constant;
    -- logger for split-operator MUX_7009_inst flow-through 
    process(IMA9_7010) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_7009_inst:flowthrough inputs: " & " BITSEL_u8_u1_7004_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_7004_wire) & " type_cast_7006_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7006_wire_constant) & " type_cast_7008_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7008_wire_constant) & " outputs:" & " IMA9_7010= "  & Convert_SLV_To_Hex_String(IMA9_7010));
      --
    end process; 
    -- flow-through select operator MUX_7009_inst
    IMA9_7010 <= type_cast_7006_wire_constant when (BITSEL_u8_u1_7004_wire(0) /=  '0') else type_cast_7008_wire_constant;
    -- logger for split-operator MUX_7019_inst flow-through 
    process(IMA10_7020) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_7019_inst:flowthrough inputs: " & " BITSEL_u8_u1_7014_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_7014_wire) & " type_cast_7016_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7016_wire_constant) & " type_cast_7018_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7018_wire_constant) & " outputs:" & " IMA10_7020= "  & Convert_SLV_To_Hex_String(IMA10_7020));
      --
    end process; 
    -- flow-through select operator MUX_7019_inst
    IMA10_7020 <= type_cast_7016_wire_constant when (BITSEL_u8_u1_7014_wire(0) /=  '0') else type_cast_7018_wire_constant;
    -- logger for split-operator MUX_7029_inst flow-through 
    process(IMA11_7030) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_7029_inst:flowthrough inputs: " & " BITSEL_u8_u1_7024_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_7024_wire) & " type_cast_7026_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7026_wire_constant) & " type_cast_7028_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7028_wire_constant) & " outputs:" & " IMA11_7030= "  & Convert_SLV_To_Hex_String(IMA11_7030));
      --
    end process; 
    -- flow-through select operator MUX_7029_inst
    IMA11_7030 <= type_cast_7026_wire_constant when (BITSEL_u8_u1_7024_wire(0) /=  '0') else type_cast_7028_wire_constant;
    -- logger for split-operator MUX_7039_inst flow-through 
    process(IMA12_7040) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_7039_inst:flowthrough inputs: " & " BITSEL_u8_u1_7034_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_7034_wire) & " type_cast_7036_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7036_wire_constant) & " type_cast_7038_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7038_wire_constant) & " outputs:" & " IMA12_7040= "  & Convert_SLV_To_Hex_String(IMA12_7040));
      --
    end process; 
    -- flow-through select operator MUX_7039_inst
    IMA12_7040 <= type_cast_7036_wire_constant when (BITSEL_u8_u1_7034_wire(0) /=  '0') else type_cast_7038_wire_constant;
    -- logger for split-operator MUX_7049_inst flow-through 
    process(IMA13_7050) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_7049_inst:flowthrough inputs: " & " BITSEL_u8_u1_7044_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_7044_wire) & " type_cast_7046_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7046_wire_constant) & " type_cast_7048_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7048_wire_constant) & " outputs:" & " IMA13_7050= "  & Convert_SLV_To_Hex_String(IMA13_7050));
      --
    end process; 
    -- flow-through select operator MUX_7049_inst
    IMA13_7050 <= type_cast_7046_wire_constant when (BITSEL_u8_u1_7044_wire(0) /=  '0') else type_cast_7048_wire_constant;
    -- logger for split-operator MUX_7059_inst flow-through 
    process(IMA14_7060) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_7059_inst:flowthrough inputs: " & " BITSEL_u8_u1_7054_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_7054_wire) & " type_cast_7056_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7056_wire_constant) & " type_cast_7058_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7058_wire_constant) & " outputs:" & " IMA14_7060= "  & Convert_SLV_To_Hex_String(IMA14_7060));
      --
    end process; 
    -- flow-through select operator MUX_7059_inst
    IMA14_7060 <= type_cast_7056_wire_constant when (BITSEL_u8_u1_7054_wire(0) /=  '0') else type_cast_7058_wire_constant;
    -- logger for split-operator MUX_7069_inst flow-through 
    process(IMA15_7070) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_7069_inst:flowthrough inputs: " & " BITSEL_u8_u1_7064_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_7064_wire) & " type_cast_7066_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7066_wire_constant) & " type_cast_7068_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7068_wire_constant) & " outputs:" & " IMA15_7070= "  & Convert_SLV_To_Hex_String(IMA15_7070));
      --
    end process; 
    -- flow-through select operator MUX_7069_inst
    IMA15_7070 <= type_cast_7066_wire_constant when (BITSEL_u8_u1_7064_wire(0) /=  '0') else type_cast_7068_wire_constant;
    -- logger for split-operator MUX_7079_inst flow-through 
    process(IMA16_7080) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_7079_inst:flowthrough inputs: " & " BITSEL_u8_u1_7074_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_7074_wire) & " type_cast_7076_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7076_wire_constant) & " type_cast_7078_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7078_wire_constant) & " outputs:" & " IMA16_7080= "  & Convert_SLV_To_Hex_String(IMA16_7080));
      --
    end process; 
    -- flow-through select operator MUX_7079_inst
    IMA16_7080 <= type_cast_7076_wire_constant when (BITSEL_u8_u1_7074_wire(0) /=  '0') else type_cast_7078_wire_constant;
    -- logger for split-operator MUX_7089_inst flow-through 
    process(IMA17_7090) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_7089_inst:flowthrough inputs: " & " BITSEL_u8_u1_7084_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_7084_wire) & " type_cast_7086_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7086_wire_constant) & " type_cast_7088_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7088_wire_constant) & " outputs:" & " IMA17_7090= "  & Convert_SLV_To_Hex_String(IMA17_7090));
      --
    end process; 
    -- flow-through select operator MUX_7089_inst
    IMA17_7090 <= type_cast_7086_wire_constant when (BITSEL_u8_u1_7084_wire(0) /=  '0') else type_cast_7088_wire_constant;
    -- logger for split-operator MUX_7099_inst flow-through 
    process(IMA18_7100) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_7099_inst:flowthrough inputs: " & " BITSEL_u8_u1_7094_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_7094_wire) & " type_cast_7096_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7096_wire_constant) & " type_cast_7098_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7098_wire_constant) & " outputs:" & " IMA18_7100= "  & Convert_SLV_To_Hex_String(IMA18_7100));
      --
    end process; 
    -- flow-through select operator MUX_7099_inst
    IMA18_7100 <= type_cast_7096_wire_constant when (BITSEL_u8_u1_7094_wire(0) /=  '0') else type_cast_7098_wire_constant;
    -- logger for split-operator MUX_7109_inst flow-through 
    process(IMA19_7110) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_7109_inst:flowthrough inputs: " & " BITSEL_u8_u1_7104_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_7104_wire) & " type_cast_7106_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7106_wire_constant) & " type_cast_7108_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7108_wire_constant) & " outputs:" & " IMA19_7110= "  & Convert_SLV_To_Hex_String(IMA19_7110));
      --
    end process; 
    -- flow-through select operator MUX_7109_inst
    IMA19_7110 <= type_cast_7106_wire_constant when (BITSEL_u8_u1_7104_wire(0) /=  '0') else type_cast_7108_wire_constant;
    -- logger for split-operator MUX_7119_inst flow-through 
    process(IMA20_7120) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_7119_inst:flowthrough inputs: " & " BITSEL_u8_u1_7114_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_7114_wire) & " type_cast_7116_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7116_wire_constant) & " type_cast_7118_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7118_wire_constant) & " outputs:" & " IMA20_7120= "  & Convert_SLV_To_Hex_String(IMA20_7120));
      --
    end process; 
    -- flow-through select operator MUX_7119_inst
    IMA20_7120 <= type_cast_7116_wire_constant when (BITSEL_u8_u1_7114_wire(0) /=  '0') else type_cast_7118_wire_constant;
    -- logger for split-operator MUX_7129_inst flow-through 
    process(IMA21_7130) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_7129_inst:flowthrough inputs: " & " BITSEL_u8_u1_7124_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_7124_wire) & " type_cast_7126_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7126_wire_constant) & " type_cast_7128_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7128_wire_constant) & " outputs:" & " IMA21_7130= "  & Convert_SLV_To_Hex_String(IMA21_7130));
      --
    end process; 
    -- flow-through select operator MUX_7129_inst
    IMA21_7130 <= type_cast_7126_wire_constant when (BITSEL_u8_u1_7124_wire(0) /=  '0') else type_cast_7128_wire_constant;
    -- logger for split-operator MUX_7139_inst flow-through 
    process(IMA22_7140) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_7139_inst:flowthrough inputs: " & " BITSEL_u8_u1_7134_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_7134_wire) & " type_cast_7136_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7136_wire_constant) & " type_cast_7138_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7138_wire_constant) & " outputs:" & " IMA22_7140= "  & Convert_SLV_To_Hex_String(IMA22_7140));
      --
    end process; 
    -- flow-through select operator MUX_7139_inst
    IMA22_7140 <= type_cast_7136_wire_constant when (BITSEL_u8_u1_7134_wire(0) /=  '0') else type_cast_7138_wire_constant;
    -- logger for split-operator MUX_7149_inst flow-through 
    process(IMA23_7150) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_7149_inst:flowthrough inputs: " & " BITSEL_u8_u1_7144_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_7144_wire) & " type_cast_7146_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7146_wire_constant) & " type_cast_7148_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7148_wire_constant) & " outputs:" & " IMA23_7150= "  & Convert_SLV_To_Hex_String(IMA23_7150));
      --
    end process; 
    -- flow-through select operator MUX_7149_inst
    IMA23_7150 <= type_cast_7146_wire_constant when (BITSEL_u8_u1_7144_wire(0) /=  '0') else type_cast_7148_wire_constant;
    -- logger for split-operator MUX_7159_inst flow-through 
    process(IMA24_7160) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_7159_inst:flowthrough inputs: " & " BITSEL_u8_u1_7154_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_7154_wire) & " type_cast_7156_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7156_wire_constant) & " type_cast_7158_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7158_wire_constant) & " outputs:" & " IMA24_7160= "  & Convert_SLV_To_Hex_String(IMA24_7160));
      --
    end process; 
    -- flow-through select operator MUX_7159_inst
    IMA24_7160 <= type_cast_7156_wire_constant when (BITSEL_u8_u1_7154_wire(0) /=  '0') else type_cast_7158_wire_constant;
    -- logger for split-operator MUX_7169_inst flow-through 
    process(IMA25_7170) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_7169_inst:flowthrough inputs: " & " BITSEL_u8_u1_7164_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_7164_wire) & " type_cast_7166_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7166_wire_constant) & " type_cast_7168_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7168_wire_constant) & " outputs:" & " IMA25_7170= "  & Convert_SLV_To_Hex_String(IMA25_7170));
      --
    end process; 
    -- flow-through select operator MUX_7169_inst
    IMA25_7170 <= type_cast_7166_wire_constant when (BITSEL_u8_u1_7164_wire(0) /=  '0') else type_cast_7168_wire_constant;
    -- logger for split-operator MUX_7179_inst flow-through 
    process(IMA26_7180) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_7179_inst:flowthrough inputs: " & " BITSEL_u8_u1_7174_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_7174_wire) & " type_cast_7176_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7176_wire_constant) & " type_cast_7178_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7178_wire_constant) & " outputs:" & " IMA26_7180= "  & Convert_SLV_To_Hex_String(IMA26_7180));
      --
    end process; 
    -- flow-through select operator MUX_7179_inst
    IMA26_7180 <= type_cast_7176_wire_constant when (BITSEL_u8_u1_7174_wire(0) /=  '0') else type_cast_7178_wire_constant;
    -- logger for split-operator MUX_7189_inst flow-through 
    process(IMA27_7190) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_7189_inst:flowthrough inputs: " & " BITSEL_u8_u1_7184_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_7184_wire) & " type_cast_7186_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7186_wire_constant) & " type_cast_7188_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7188_wire_constant) & " outputs:" & " IMA27_7190= "  & Convert_SLV_To_Hex_String(IMA27_7190));
      --
    end process; 
    -- flow-through select operator MUX_7189_inst
    IMA27_7190 <= type_cast_7186_wire_constant when (BITSEL_u8_u1_7184_wire(0) /=  '0') else type_cast_7188_wire_constant;
    -- logger for split-operator MUX_7199_inst flow-through 
    process(IMA28_7200) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_7199_inst:flowthrough inputs: " & " BITSEL_u8_u1_7194_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_7194_wire) & " type_cast_7196_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7196_wire_constant) & " type_cast_7198_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7198_wire_constant) & " outputs:" & " IMA28_7200= "  & Convert_SLV_To_Hex_String(IMA28_7200));
      --
    end process; 
    -- flow-through select operator MUX_7199_inst
    IMA28_7200 <= type_cast_7196_wire_constant when (BITSEL_u8_u1_7194_wire(0) /=  '0') else type_cast_7198_wire_constant;
    -- logger for split-operator MUX_7209_inst flow-through 
    process(IMA29_7210) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_7209_inst:flowthrough inputs: " & " BITSEL_u8_u1_7204_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_7204_wire) & " type_cast_7206_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7206_wire_constant) & " type_cast_7208_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7208_wire_constant) & " outputs:" & " IMA29_7210= "  & Convert_SLV_To_Hex_String(IMA29_7210));
      --
    end process; 
    -- flow-through select operator MUX_7209_inst
    IMA29_7210 <= type_cast_7206_wire_constant when (BITSEL_u8_u1_7204_wire(0) /=  '0') else type_cast_7208_wire_constant;
    -- logger for split-operator MUX_7219_inst flow-through 
    process(IMA30_7220) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_7219_inst:flowthrough inputs: " & " BITSEL_u8_u1_7214_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_7214_wire) & " type_cast_7216_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7216_wire_constant) & " type_cast_7218_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7218_wire_constant) & " outputs:" & " IMA30_7220= "  & Convert_SLV_To_Hex_String(IMA30_7220));
      --
    end process; 
    -- flow-through select operator MUX_7219_inst
    IMA30_7220 <= type_cast_7216_wire_constant when (BITSEL_u8_u1_7214_wire(0) /=  '0') else type_cast_7218_wire_constant;
    -- logger for split-operator MUX_7229_inst flow-through 
    process(IMA31_7230) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_7229_inst:flowthrough inputs: " & " BITSEL_u8_u1_7224_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_7224_wire) & " type_cast_7226_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7226_wire_constant) & " type_cast_7228_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7228_wire_constant) & " outputs:" & " IMA31_7230= "  & Convert_SLV_To_Hex_String(IMA31_7230));
      --
    end process; 
    -- flow-through select operator MUX_7229_inst
    IMA31_7230 <= type_cast_7226_wire_constant when (BITSEL_u8_u1_7224_wire(0) /=  '0') else type_cast_7228_wire_constant;
    -- logger for split-operator MUX_7239_inst flow-through 
    process(IMA32_7240) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_7239_inst:flowthrough inputs: " & " BITSEL_u8_u1_7234_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_7234_wire) & " type_cast_7236_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7236_wire_constant) & " type_cast_7238_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7238_wire_constant) & " outputs:" & " IMA32_7240= "  & Convert_SLV_To_Hex_String(IMA32_7240));
      --
    end process; 
    -- flow-through select operator MUX_7239_inst
    IMA32_7240 <= type_cast_7236_wire_constant when (BITSEL_u8_u1_7234_wire(0) /=  '0') else type_cast_7238_wire_constant;
    -- logger for split-operator MUX_7249_inst flow-through 
    process(IMA33_7250) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_7249_inst:flowthrough inputs: " & " BITSEL_u8_u1_7244_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_7244_wire) & " type_cast_7246_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7246_wire_constant) & " type_cast_7248_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7248_wire_constant) & " outputs:" & " IMA33_7250= "  & Convert_SLV_To_Hex_String(IMA33_7250));
      --
    end process; 
    -- flow-through select operator MUX_7249_inst
    IMA33_7250 <= type_cast_7246_wire_constant when (BITSEL_u8_u1_7244_wire(0) /=  '0') else type_cast_7248_wire_constant;
    -- logger for split-operator MUX_7259_inst flow-through 
    process(IMA34_7260) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_7259_inst:flowthrough inputs: " & " BITSEL_u8_u1_7254_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_7254_wire) & " type_cast_7256_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7256_wire_constant) & " type_cast_7258_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7258_wire_constant) & " outputs:" & " IMA34_7260= "  & Convert_SLV_To_Hex_String(IMA34_7260));
      --
    end process; 
    -- flow-through select operator MUX_7259_inst
    IMA34_7260 <= type_cast_7256_wire_constant when (BITSEL_u8_u1_7254_wire(0) /=  '0') else type_cast_7258_wire_constant;
    -- logger for split-operator MUX_7269_inst flow-through 
    process(IMA35_7270) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_7269_inst:flowthrough inputs: " & " BITSEL_u8_u1_7264_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_7264_wire) & " type_cast_7266_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7266_wire_constant) & " type_cast_7268_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7268_wire_constant) & " outputs:" & " IMA35_7270= "  & Convert_SLV_To_Hex_String(IMA35_7270));
      --
    end process; 
    -- flow-through select operator MUX_7269_inst
    IMA35_7270 <= type_cast_7266_wire_constant when (BITSEL_u8_u1_7264_wire(0) /=  '0') else type_cast_7268_wire_constant;
    -- logger for split-operator MUX_7279_inst flow-through 
    process(IMA36_7280) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_7279_inst:flowthrough inputs: " & " BITSEL_u8_u1_7274_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_7274_wire) & " type_cast_7276_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7276_wire_constant) & " type_cast_7278_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7278_wire_constant) & " outputs:" & " IMA36_7280= "  & Convert_SLV_To_Hex_String(IMA36_7280));
      --
    end process; 
    -- flow-through select operator MUX_7279_inst
    IMA36_7280 <= type_cast_7276_wire_constant when (BITSEL_u8_u1_7274_wire(0) /=  '0') else type_cast_7278_wire_constant;
    -- logger for split-operator MUX_7289_inst flow-through 
    process(IMA37_7290) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_7289_inst:flowthrough inputs: " & " BITSEL_u8_u1_7284_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_7284_wire) & " type_cast_7286_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7286_wire_constant) & " type_cast_7288_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7288_wire_constant) & " outputs:" & " IMA37_7290= "  & Convert_SLV_To_Hex_String(IMA37_7290));
      --
    end process; 
    -- flow-through select operator MUX_7289_inst
    IMA37_7290 <= type_cast_7286_wire_constant when (BITSEL_u8_u1_7284_wire(0) /=  '0') else type_cast_7288_wire_constant;
    -- logger for split-operator MUX_7299_inst flow-through 
    process(IMA38_7300) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_7299_inst:flowthrough inputs: " & " BITSEL_u8_u1_7294_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_7294_wire) & " type_cast_7296_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7296_wire_constant) & " type_cast_7298_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7298_wire_constant) & " outputs:" & " IMA38_7300= "  & Convert_SLV_To_Hex_String(IMA38_7300));
      --
    end process; 
    -- flow-through select operator MUX_7299_inst
    IMA38_7300 <= type_cast_7296_wire_constant when (BITSEL_u8_u1_7294_wire(0) /=  '0') else type_cast_7298_wire_constant;
    -- logger for split-operator MUX_7309_inst flow-through 
    process(IMA39_7310) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_7309_inst:flowthrough inputs: " & " BITSEL_u8_u1_7304_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_7304_wire) & " type_cast_7306_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7306_wire_constant) & " type_cast_7308_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7308_wire_constant) & " outputs:" & " IMA39_7310= "  & Convert_SLV_To_Hex_String(IMA39_7310));
      --
    end process; 
    -- flow-through select operator MUX_7309_inst
    IMA39_7310 <= type_cast_7306_wire_constant when (BITSEL_u8_u1_7304_wire(0) /=  '0') else type_cast_7308_wire_constant;
    -- logger for split-operator MUX_7319_inst flow-through 
    process(IMA40_7320) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_7319_inst:flowthrough inputs: " & " BITSEL_u8_u1_7314_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_7314_wire) & " type_cast_7316_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7316_wire_constant) & " type_cast_7318_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7318_wire_constant) & " outputs:" & " IMA40_7320= "  & Convert_SLV_To_Hex_String(IMA40_7320));
      --
    end process; 
    -- flow-through select operator MUX_7319_inst
    IMA40_7320 <= type_cast_7316_wire_constant when (BITSEL_u8_u1_7314_wire(0) /=  '0') else type_cast_7318_wire_constant;
    -- logger for split-operator MUX_7329_inst flow-through 
    process(IMA41_7330) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_7329_inst:flowthrough inputs: " & " BITSEL_u8_u1_7324_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_7324_wire) & " type_cast_7326_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7326_wire_constant) & " type_cast_7328_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7328_wire_constant) & " outputs:" & " IMA41_7330= "  & Convert_SLV_To_Hex_String(IMA41_7330));
      --
    end process; 
    -- flow-through select operator MUX_7329_inst
    IMA41_7330 <= type_cast_7326_wire_constant when (BITSEL_u8_u1_7324_wire(0) /=  '0') else type_cast_7328_wire_constant;
    -- logger for split-operator MUX_7339_inst flow-through 
    process(IMA42_7340) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_7339_inst:flowthrough inputs: " & " BITSEL_u8_u1_7334_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_7334_wire) & " type_cast_7336_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7336_wire_constant) & " type_cast_7338_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7338_wire_constant) & " outputs:" & " IMA42_7340= "  & Convert_SLV_To_Hex_String(IMA42_7340));
      --
    end process; 
    -- flow-through select operator MUX_7339_inst
    IMA42_7340 <= type_cast_7336_wire_constant when (BITSEL_u8_u1_7334_wire(0) /=  '0') else type_cast_7338_wire_constant;
    -- logger for split-operator MUX_7349_inst flow-through 
    process(IMA43_7350) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_7349_inst:flowthrough inputs: " & " BITSEL_u8_u1_7344_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_7344_wire) & " type_cast_7346_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7346_wire_constant) & " type_cast_7348_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7348_wire_constant) & " outputs:" & " IMA43_7350= "  & Convert_SLV_To_Hex_String(IMA43_7350));
      --
    end process; 
    -- flow-through select operator MUX_7349_inst
    IMA43_7350 <= type_cast_7346_wire_constant when (BITSEL_u8_u1_7344_wire(0) /=  '0') else type_cast_7348_wire_constant;
    -- logger for split-operator MUX_7359_inst flow-through 
    process(IMA44_7360) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_7359_inst:flowthrough inputs: " & " BITSEL_u8_u1_7354_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_7354_wire) & " type_cast_7356_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7356_wire_constant) & " type_cast_7358_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7358_wire_constant) & " outputs:" & " IMA44_7360= "  & Convert_SLV_To_Hex_String(IMA44_7360));
      --
    end process; 
    -- flow-through select operator MUX_7359_inst
    IMA44_7360 <= type_cast_7356_wire_constant when (BITSEL_u8_u1_7354_wire(0) /=  '0') else type_cast_7358_wire_constant;
    -- logger for split-operator MUX_7369_inst flow-through 
    process(IMA45_7370) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_7369_inst:flowthrough inputs: " & " BITSEL_u8_u1_7364_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_7364_wire) & " type_cast_7366_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7366_wire_constant) & " type_cast_7368_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7368_wire_constant) & " outputs:" & " IMA45_7370= "  & Convert_SLV_To_Hex_String(IMA45_7370));
      --
    end process; 
    -- flow-through select operator MUX_7369_inst
    IMA45_7370 <= type_cast_7366_wire_constant when (BITSEL_u8_u1_7364_wire(0) /=  '0') else type_cast_7368_wire_constant;
    -- logger for split-operator MUX_7379_inst flow-through 
    process(IMA46_7380) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_7379_inst:flowthrough inputs: " & " BITSEL_u8_u1_7374_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_7374_wire) & " type_cast_7376_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7376_wire_constant) & " type_cast_7378_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7378_wire_constant) & " outputs:" & " IMA46_7380= "  & Convert_SLV_To_Hex_String(IMA46_7380));
      --
    end process; 
    -- flow-through select operator MUX_7379_inst
    IMA46_7380 <= type_cast_7376_wire_constant when (BITSEL_u8_u1_7374_wire(0) /=  '0') else type_cast_7378_wire_constant;
    -- logger for split-operator MUX_7389_inst flow-through 
    process(IMA47_7390) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_7389_inst:flowthrough inputs: " & " BITSEL_u8_u1_7384_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_7384_wire) & " type_cast_7386_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7386_wire_constant) & " type_cast_7388_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7388_wire_constant) & " outputs:" & " IMA47_7390= "  & Convert_SLV_To_Hex_String(IMA47_7390));
      --
    end process; 
    -- flow-through select operator MUX_7389_inst
    IMA47_7390 <= type_cast_7386_wire_constant when (BITSEL_u8_u1_7384_wire(0) /=  '0') else type_cast_7388_wire_constant;
    -- logger for split-operator MUX_7399_inst flow-through 
    process(IMA48_7400) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_7399_inst:flowthrough inputs: " & " BITSEL_u8_u1_7394_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_7394_wire) & " type_cast_7396_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7396_wire_constant) & " type_cast_7398_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7398_wire_constant) & " outputs:" & " IMA48_7400= "  & Convert_SLV_To_Hex_String(IMA48_7400));
      --
    end process; 
    -- flow-through select operator MUX_7399_inst
    IMA48_7400 <= type_cast_7396_wire_constant when (BITSEL_u8_u1_7394_wire(0) /=  '0') else type_cast_7398_wire_constant;
    -- logger for split-operator MUX_7409_inst flow-through 
    process(IMA49_7410) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_7409_inst:flowthrough inputs: " & " BITSEL_u8_u1_7404_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_7404_wire) & " type_cast_7406_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7406_wire_constant) & " type_cast_7408_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7408_wire_constant) & " outputs:" & " IMA49_7410= "  & Convert_SLV_To_Hex_String(IMA49_7410));
      --
    end process; 
    -- flow-through select operator MUX_7409_inst
    IMA49_7410 <= type_cast_7406_wire_constant when (BITSEL_u8_u1_7404_wire(0) /=  '0') else type_cast_7408_wire_constant;
    -- logger for split-operator MUX_7419_inst flow-through 
    process(IMA50_7420) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_7419_inst:flowthrough inputs: " & " BITSEL_u8_u1_7414_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_7414_wire) & " type_cast_7416_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7416_wire_constant) & " type_cast_7418_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7418_wire_constant) & " outputs:" & " IMA50_7420= "  & Convert_SLV_To_Hex_String(IMA50_7420));
      --
    end process; 
    -- flow-through select operator MUX_7419_inst
    IMA50_7420 <= type_cast_7416_wire_constant when (BITSEL_u8_u1_7414_wire(0) /=  '0') else type_cast_7418_wire_constant;
    -- logger for split-operator MUX_7429_inst flow-through 
    process(IMA51_7430) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_7429_inst:flowthrough inputs: " & " BITSEL_u8_u1_7424_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_7424_wire) & " type_cast_7426_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7426_wire_constant) & " type_cast_7428_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7428_wire_constant) & " outputs:" & " IMA51_7430= "  & Convert_SLV_To_Hex_String(IMA51_7430));
      --
    end process; 
    -- flow-through select operator MUX_7429_inst
    IMA51_7430 <= type_cast_7426_wire_constant when (BITSEL_u8_u1_7424_wire(0) /=  '0') else type_cast_7428_wire_constant;
    -- logger for split-operator MUX_7439_inst flow-through 
    process(IMA52_7440) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_7439_inst:flowthrough inputs: " & " BITSEL_u8_u1_7434_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_7434_wire) & " type_cast_7436_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7436_wire_constant) & " type_cast_7438_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7438_wire_constant) & " outputs:" & " IMA52_7440= "  & Convert_SLV_To_Hex_String(IMA52_7440));
      --
    end process; 
    -- flow-through select operator MUX_7439_inst
    IMA52_7440 <= type_cast_7436_wire_constant when (BITSEL_u8_u1_7434_wire(0) /=  '0') else type_cast_7438_wire_constant;
    -- logger for split-operator MUX_7449_inst flow-through 
    process(IMA53_7450) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_7449_inst:flowthrough inputs: " & " BITSEL_u8_u1_7444_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_7444_wire) & " type_cast_7446_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7446_wire_constant) & " type_cast_7448_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7448_wire_constant) & " outputs:" & " IMA53_7450= "  & Convert_SLV_To_Hex_String(IMA53_7450));
      --
    end process; 
    -- flow-through select operator MUX_7449_inst
    IMA53_7450 <= type_cast_7446_wire_constant when (BITSEL_u8_u1_7444_wire(0) /=  '0') else type_cast_7448_wire_constant;
    -- logger for split-operator MUX_7459_inst flow-through 
    process(IMA54_7460) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_7459_inst:flowthrough inputs: " & " BITSEL_u8_u1_7454_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_7454_wire) & " type_cast_7456_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7456_wire_constant) & " type_cast_7458_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7458_wire_constant) & " outputs:" & " IMA54_7460= "  & Convert_SLV_To_Hex_String(IMA54_7460));
      --
    end process; 
    -- flow-through select operator MUX_7459_inst
    IMA54_7460 <= type_cast_7456_wire_constant when (BITSEL_u8_u1_7454_wire(0) /=  '0') else type_cast_7458_wire_constant;
    -- logger for split-operator MUX_7469_inst flow-through 
    process(IMA55_7470) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_7469_inst:flowthrough inputs: " & " BITSEL_u8_u1_7464_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_7464_wire) & " type_cast_7466_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7466_wire_constant) & " type_cast_7468_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7468_wire_constant) & " outputs:" & " IMA55_7470= "  & Convert_SLV_To_Hex_String(IMA55_7470));
      --
    end process; 
    -- flow-through select operator MUX_7469_inst
    IMA55_7470 <= type_cast_7466_wire_constant when (BITSEL_u8_u1_7464_wire(0) /=  '0') else type_cast_7468_wire_constant;
    -- logger for split-operator MUX_7479_inst flow-through 
    process(IMA56_7480) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_7479_inst:flowthrough inputs: " & " BITSEL_u8_u1_7474_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_7474_wire) & " type_cast_7476_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7476_wire_constant) & " type_cast_7478_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7478_wire_constant) & " outputs:" & " IMA56_7480= "  & Convert_SLV_To_Hex_String(IMA56_7480));
      --
    end process; 
    -- flow-through select operator MUX_7479_inst
    IMA56_7480 <= type_cast_7476_wire_constant when (BITSEL_u8_u1_7474_wire(0) /=  '0') else type_cast_7478_wire_constant;
    -- logger for split-operator MUX_7489_inst flow-through 
    process(IMA57_7490) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_7489_inst:flowthrough inputs: " & " BITSEL_u8_u1_7484_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_7484_wire) & " type_cast_7486_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7486_wire_constant) & " type_cast_7488_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7488_wire_constant) & " outputs:" & " IMA57_7490= "  & Convert_SLV_To_Hex_String(IMA57_7490));
      --
    end process; 
    -- flow-through select operator MUX_7489_inst
    IMA57_7490 <= type_cast_7486_wire_constant when (BITSEL_u8_u1_7484_wire(0) /=  '0') else type_cast_7488_wire_constant;
    -- logger for split-operator MUX_7499_inst flow-through 
    process(IMA58_7500) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_7499_inst:flowthrough inputs: " & " BITSEL_u8_u1_7494_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_7494_wire) & " type_cast_7496_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7496_wire_constant) & " type_cast_7498_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7498_wire_constant) & " outputs:" & " IMA58_7500= "  & Convert_SLV_To_Hex_String(IMA58_7500));
      --
    end process; 
    -- flow-through select operator MUX_7499_inst
    IMA58_7500 <= type_cast_7496_wire_constant when (BITSEL_u8_u1_7494_wire(0) /=  '0') else type_cast_7498_wire_constant;
    -- logger for split-operator MUX_7509_inst flow-through 
    process(IMA59_7510) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_7509_inst:flowthrough inputs: " & " BITSEL_u8_u1_7504_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_7504_wire) & " type_cast_7506_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7506_wire_constant) & " type_cast_7508_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7508_wire_constant) & " outputs:" & " IMA59_7510= "  & Convert_SLV_To_Hex_String(IMA59_7510));
      --
    end process; 
    -- flow-through select operator MUX_7509_inst
    IMA59_7510 <= type_cast_7506_wire_constant when (BITSEL_u8_u1_7504_wire(0) /=  '0') else type_cast_7508_wire_constant;
    -- logger for split-operator MUX_7519_inst flow-through 
    process(IMA60_7520) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_7519_inst:flowthrough inputs: " & " BITSEL_u8_u1_7514_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_7514_wire) & " type_cast_7516_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7516_wire_constant) & " type_cast_7518_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7518_wire_constant) & " outputs:" & " IMA60_7520= "  & Convert_SLV_To_Hex_String(IMA60_7520));
      --
    end process; 
    -- flow-through select operator MUX_7519_inst
    IMA60_7520 <= type_cast_7516_wire_constant when (BITSEL_u8_u1_7514_wire(0) /=  '0') else type_cast_7518_wire_constant;
    -- logger for split-operator MUX_7529_inst flow-through 
    process(IMA61_7530) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_7529_inst:flowthrough inputs: " & " BITSEL_u8_u1_7524_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_7524_wire) & " type_cast_7526_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7526_wire_constant) & " type_cast_7528_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7528_wire_constant) & " outputs:" & " IMA61_7530= "  & Convert_SLV_To_Hex_String(IMA61_7530));
      --
    end process; 
    -- flow-through select operator MUX_7529_inst
    IMA61_7530 <= type_cast_7526_wire_constant when (BITSEL_u8_u1_7524_wire(0) /=  '0') else type_cast_7528_wire_constant;
    -- logger for split-operator MUX_7539_inst flow-through 
    process(IMA62_7540) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_7539_inst:flowthrough inputs: " & " BITSEL_u8_u1_7534_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_7534_wire) & " type_cast_7536_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7536_wire_constant) & " type_cast_7538_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7538_wire_constant) & " outputs:" & " IMA62_7540= "  & Convert_SLV_To_Hex_String(IMA62_7540));
      --
    end process; 
    -- flow-through select operator MUX_7539_inst
    IMA62_7540 <= type_cast_7536_wire_constant when (BITSEL_u8_u1_7534_wire(0) /=  '0') else type_cast_7538_wire_constant;
    -- logger for split-operator MUX_7549_inst flow-through 
    process(IMA63_7550) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_7549_inst:flowthrough inputs: " & " BITSEL_u8_u1_7544_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_7544_wire) & " type_cast_7546_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7546_wire_constant) & " type_cast_7548_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7548_wire_constant) & " outputs:" & " IMA63_7550= "  & Convert_SLV_To_Hex_String(IMA63_7550));
      --
    end process; 
    -- flow-through select operator MUX_7549_inst
    IMA63_7550 <= type_cast_7546_wire_constant when (BITSEL_u8_u1_7544_wire(0) /=  '0') else type_cast_7548_wire_constant;
    -- logger for split-operator MUX_7559_inst flow-through 
    process(IMA64_7560) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_7559_inst:flowthrough inputs: " & " BITSEL_u8_u1_7554_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_7554_wire) & " type_cast_7556_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7556_wire_constant) & " type_cast_7558_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7558_wire_constant) & " outputs:" & " IMA64_7560= "  & Convert_SLV_To_Hex_String(IMA64_7560));
      --
    end process; 
    -- flow-through select operator MUX_7559_inst
    IMA64_7560 <= type_cast_7556_wire_constant when (BITSEL_u8_u1_7554_wire(0) /=  '0') else type_cast_7558_wire_constant;
    -- logger for split-operator MUX_7569_inst flow-through 
    process(IMA65_7570) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_7569_inst:flowthrough inputs: " & " BITSEL_u8_u1_7564_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_7564_wire) & " type_cast_7566_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7566_wire_constant) & " type_cast_7568_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7568_wire_constant) & " outputs:" & " IMA65_7570= "  & Convert_SLV_To_Hex_String(IMA65_7570));
      --
    end process; 
    -- flow-through select operator MUX_7569_inst
    IMA65_7570 <= type_cast_7566_wire_constant when (BITSEL_u8_u1_7564_wire(0) /=  '0') else type_cast_7568_wire_constant;
    -- logger for split-operator MUX_7579_inst flow-through 
    process(IMA66_7580) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_7579_inst:flowthrough inputs: " & " BITSEL_u8_u1_7574_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_7574_wire) & " type_cast_7576_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7576_wire_constant) & " type_cast_7578_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7578_wire_constant) & " outputs:" & " IMA66_7580= "  & Convert_SLV_To_Hex_String(IMA66_7580));
      --
    end process; 
    -- flow-through select operator MUX_7579_inst
    IMA66_7580 <= type_cast_7576_wire_constant when (BITSEL_u8_u1_7574_wire(0) /=  '0') else type_cast_7578_wire_constant;
    -- logger for split-operator MUX_7589_inst flow-through 
    process(IMA67_7590) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_7589_inst:flowthrough inputs: " & " BITSEL_u8_u1_7584_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_7584_wire) & " type_cast_7586_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7586_wire_constant) & " type_cast_7588_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7588_wire_constant) & " outputs:" & " IMA67_7590= "  & Convert_SLV_To_Hex_String(IMA67_7590));
      --
    end process; 
    -- flow-through select operator MUX_7589_inst
    IMA67_7590 <= type_cast_7586_wire_constant when (BITSEL_u8_u1_7584_wire(0) /=  '0') else type_cast_7588_wire_constant;
    -- logger for split-operator MUX_7599_inst flow-through 
    process(IMA68_7600) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_7599_inst:flowthrough inputs: " & " BITSEL_u8_u1_7594_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_7594_wire) & " type_cast_7596_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7596_wire_constant) & " type_cast_7598_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7598_wire_constant) & " outputs:" & " IMA68_7600= "  & Convert_SLV_To_Hex_String(IMA68_7600));
      --
    end process; 
    -- flow-through select operator MUX_7599_inst
    IMA68_7600 <= type_cast_7596_wire_constant when (BITSEL_u8_u1_7594_wire(0) /=  '0') else type_cast_7598_wire_constant;
    -- logger for split-operator MUX_7609_inst flow-through 
    process(IMA69_7610) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_7609_inst:flowthrough inputs: " & " BITSEL_u8_u1_7604_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_7604_wire) & " type_cast_7606_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7606_wire_constant) & " type_cast_7608_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7608_wire_constant) & " outputs:" & " IMA69_7610= "  & Convert_SLV_To_Hex_String(IMA69_7610));
      --
    end process; 
    -- flow-through select operator MUX_7609_inst
    IMA69_7610 <= type_cast_7606_wire_constant when (BITSEL_u8_u1_7604_wire(0) /=  '0') else type_cast_7608_wire_constant;
    -- logger for split-operator MUX_7619_inst flow-through 
    process(IMA70_7620) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_7619_inst:flowthrough inputs: " & " BITSEL_u8_u1_7614_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_7614_wire) & " type_cast_7616_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7616_wire_constant) & " type_cast_7618_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7618_wire_constant) & " outputs:" & " IMA70_7620= "  & Convert_SLV_To_Hex_String(IMA70_7620));
      --
    end process; 
    -- flow-through select operator MUX_7619_inst
    IMA70_7620 <= type_cast_7616_wire_constant when (BITSEL_u8_u1_7614_wire(0) /=  '0') else type_cast_7618_wire_constant;
    -- logger for split-operator MUX_7629_inst flow-through 
    process(IMA71_7630) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_7629_inst:flowthrough inputs: " & " BITSEL_u8_u1_7624_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_7624_wire) & " type_cast_7626_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7626_wire_constant) & " type_cast_7628_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7628_wire_constant) & " outputs:" & " IMA71_7630= "  & Convert_SLV_To_Hex_String(IMA71_7630));
      --
    end process; 
    -- flow-through select operator MUX_7629_inst
    IMA71_7630 <= type_cast_7626_wire_constant when (BITSEL_u8_u1_7624_wire(0) /=  '0') else type_cast_7628_wire_constant;
    -- logger for split-operator MUX_7639_inst flow-through 
    process(IMA72_7640) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_7639_inst:flowthrough inputs: " & " BITSEL_u8_u1_7634_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_7634_wire) & " type_cast_7636_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7636_wire_constant) & " type_cast_7638_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7638_wire_constant) & " outputs:" & " IMA72_7640= "  & Convert_SLV_To_Hex_String(IMA72_7640));
      --
    end process; 
    -- flow-through select operator MUX_7639_inst
    IMA72_7640 <= type_cast_7636_wire_constant when (BITSEL_u8_u1_7634_wire(0) /=  '0') else type_cast_7638_wire_constant;
    -- logger for split-operator MUX_7649_inst flow-through 
    process(IMA73_7650) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_7649_inst:flowthrough inputs: " & " BITSEL_u8_u1_7644_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_7644_wire) & " type_cast_7646_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7646_wire_constant) & " type_cast_7648_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7648_wire_constant) & " outputs:" & " IMA73_7650= "  & Convert_SLV_To_Hex_String(IMA73_7650));
      --
    end process; 
    -- flow-through select operator MUX_7649_inst
    IMA73_7650 <= type_cast_7646_wire_constant when (BITSEL_u8_u1_7644_wire(0) /=  '0') else type_cast_7648_wire_constant;
    -- logger for split-operator MUX_7659_inst flow-through 
    process(IMA74_7660) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_7659_inst:flowthrough inputs: " & " BITSEL_u8_u1_7654_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_7654_wire) & " type_cast_7656_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7656_wire_constant) & " type_cast_7658_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7658_wire_constant) & " outputs:" & " IMA74_7660= "  & Convert_SLV_To_Hex_String(IMA74_7660));
      --
    end process; 
    -- flow-through select operator MUX_7659_inst
    IMA74_7660 <= type_cast_7656_wire_constant when (BITSEL_u8_u1_7654_wire(0) /=  '0') else type_cast_7658_wire_constant;
    -- logger for split-operator MUX_7669_inst flow-through 
    process(IMA75_7670) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_7669_inst:flowthrough inputs: " & " BITSEL_u8_u1_7664_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_7664_wire) & " type_cast_7666_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7666_wire_constant) & " type_cast_7668_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7668_wire_constant) & " outputs:" & " IMA75_7670= "  & Convert_SLV_To_Hex_String(IMA75_7670));
      --
    end process; 
    -- flow-through select operator MUX_7669_inst
    IMA75_7670 <= type_cast_7666_wire_constant when (BITSEL_u8_u1_7664_wire(0) /=  '0') else type_cast_7668_wire_constant;
    -- logger for split-operator MUX_7679_inst flow-through 
    process(IMA76_7680) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_7679_inst:flowthrough inputs: " & " BITSEL_u8_u1_7674_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_7674_wire) & " type_cast_7676_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7676_wire_constant) & " type_cast_7678_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7678_wire_constant) & " outputs:" & " IMA76_7680= "  & Convert_SLV_To_Hex_String(IMA76_7680));
      --
    end process; 
    -- flow-through select operator MUX_7679_inst
    IMA76_7680 <= type_cast_7676_wire_constant when (BITSEL_u8_u1_7674_wire(0) /=  '0') else type_cast_7678_wire_constant;
    -- logger for split-operator MUX_7689_inst flow-through 
    process(IMA77_7690) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_7689_inst:flowthrough inputs: " & " BITSEL_u8_u1_7684_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_7684_wire) & " type_cast_7686_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7686_wire_constant) & " type_cast_7688_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7688_wire_constant) & " outputs:" & " IMA77_7690= "  & Convert_SLV_To_Hex_String(IMA77_7690));
      --
    end process; 
    -- flow-through select operator MUX_7689_inst
    IMA77_7690 <= type_cast_7686_wire_constant when (BITSEL_u8_u1_7684_wire(0) /=  '0') else type_cast_7688_wire_constant;
    -- logger for split-operator MUX_7699_inst flow-through 
    process(IMA78_7700) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_7699_inst:flowthrough inputs: " & " BITSEL_u8_u1_7694_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_7694_wire) & " type_cast_7696_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7696_wire_constant) & " type_cast_7698_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7698_wire_constant) & " outputs:" & " IMA78_7700= "  & Convert_SLV_To_Hex_String(IMA78_7700));
      --
    end process; 
    -- flow-through select operator MUX_7699_inst
    IMA78_7700 <= type_cast_7696_wire_constant when (BITSEL_u8_u1_7694_wire(0) /=  '0') else type_cast_7698_wire_constant;
    -- logger for split-operator MUX_7709_inst flow-through 
    process(IMA79_7710) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_7709_inst:flowthrough inputs: " & " BITSEL_u8_u1_7704_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_7704_wire) & " type_cast_7706_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7706_wire_constant) & " type_cast_7708_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7708_wire_constant) & " outputs:" & " IMA79_7710= "  & Convert_SLV_To_Hex_String(IMA79_7710));
      --
    end process; 
    -- flow-through select operator MUX_7709_inst
    IMA79_7710 <= type_cast_7706_wire_constant when (BITSEL_u8_u1_7704_wire(0) /=  '0') else type_cast_7708_wire_constant;
    -- logger for split-operator MUX_7719_inst flow-through 
    process(IMA80_7720) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_7719_inst:flowthrough inputs: " & " BITSEL_u8_u1_7714_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_7714_wire) & " type_cast_7716_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7716_wire_constant) & " type_cast_7718_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7718_wire_constant) & " outputs:" & " IMA80_7720= "  & Convert_SLV_To_Hex_String(IMA80_7720));
      --
    end process; 
    -- flow-through select operator MUX_7719_inst
    IMA80_7720 <= type_cast_7716_wire_constant when (BITSEL_u8_u1_7714_wire(0) /=  '0') else type_cast_7718_wire_constant;
    -- logger for split-operator MUX_7729_inst flow-through 
    process(IMA81_7730) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_7729_inst:flowthrough inputs: " & " BITSEL_u8_u1_7724_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_7724_wire) & " type_cast_7726_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7726_wire_constant) & " type_cast_7728_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7728_wire_constant) & " outputs:" & " IMA81_7730= "  & Convert_SLV_To_Hex_String(IMA81_7730));
      --
    end process; 
    -- flow-through select operator MUX_7729_inst
    IMA81_7730 <= type_cast_7726_wire_constant when (BITSEL_u8_u1_7724_wire(0) /=  '0') else type_cast_7728_wire_constant;
    -- logger for split-operator MUX_7739_inst flow-through 
    process(IMA82_7740) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_7739_inst:flowthrough inputs: " & " BITSEL_u8_u1_7734_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_7734_wire) & " type_cast_7736_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7736_wire_constant) & " type_cast_7738_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7738_wire_constant) & " outputs:" & " IMA82_7740= "  & Convert_SLV_To_Hex_String(IMA82_7740));
      --
    end process; 
    -- flow-through select operator MUX_7739_inst
    IMA82_7740 <= type_cast_7736_wire_constant when (BITSEL_u8_u1_7734_wire(0) /=  '0') else type_cast_7738_wire_constant;
    -- logger for split-operator MUX_7749_inst flow-through 
    process(IMA83_7750) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_7749_inst:flowthrough inputs: " & " BITSEL_u8_u1_7744_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_7744_wire) & " type_cast_7746_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7746_wire_constant) & " type_cast_7748_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7748_wire_constant) & " outputs:" & " IMA83_7750= "  & Convert_SLV_To_Hex_String(IMA83_7750));
      --
    end process; 
    -- flow-through select operator MUX_7749_inst
    IMA83_7750 <= type_cast_7746_wire_constant when (BITSEL_u8_u1_7744_wire(0) /=  '0') else type_cast_7748_wire_constant;
    -- logger for split-operator MUX_7759_inst flow-through 
    process(IMA84_7760) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_7759_inst:flowthrough inputs: " & " BITSEL_u8_u1_7754_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_7754_wire) & " type_cast_7756_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7756_wire_constant) & " type_cast_7758_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7758_wire_constant) & " outputs:" & " IMA84_7760= "  & Convert_SLV_To_Hex_String(IMA84_7760));
      --
    end process; 
    -- flow-through select operator MUX_7759_inst
    IMA84_7760 <= type_cast_7756_wire_constant when (BITSEL_u8_u1_7754_wire(0) /=  '0') else type_cast_7758_wire_constant;
    -- logger for split-operator MUX_7769_inst flow-through 
    process(IMA85_7770) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_7769_inst:flowthrough inputs: " & " BITSEL_u8_u1_7764_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_7764_wire) & " type_cast_7766_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7766_wire_constant) & " type_cast_7768_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7768_wire_constant) & " outputs:" & " IMA85_7770= "  & Convert_SLV_To_Hex_String(IMA85_7770));
      --
    end process; 
    -- flow-through select operator MUX_7769_inst
    IMA85_7770 <= type_cast_7766_wire_constant when (BITSEL_u8_u1_7764_wire(0) /=  '0') else type_cast_7768_wire_constant;
    -- logger for split-operator MUX_7779_inst flow-through 
    process(IMA86_7780) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_7779_inst:flowthrough inputs: " & " BITSEL_u8_u1_7774_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_7774_wire) & " type_cast_7776_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7776_wire_constant) & " type_cast_7778_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7778_wire_constant) & " outputs:" & " IMA86_7780= "  & Convert_SLV_To_Hex_String(IMA86_7780));
      --
    end process; 
    -- flow-through select operator MUX_7779_inst
    IMA86_7780 <= type_cast_7776_wire_constant when (BITSEL_u8_u1_7774_wire(0) /=  '0') else type_cast_7778_wire_constant;
    -- logger for split-operator MUX_7789_inst flow-through 
    process(IMA87_7790) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_7789_inst:flowthrough inputs: " & " BITSEL_u8_u1_7784_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_7784_wire) & " type_cast_7786_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7786_wire_constant) & " type_cast_7788_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7788_wire_constant) & " outputs:" & " IMA87_7790= "  & Convert_SLV_To_Hex_String(IMA87_7790));
      --
    end process; 
    -- flow-through select operator MUX_7789_inst
    IMA87_7790 <= type_cast_7786_wire_constant when (BITSEL_u8_u1_7784_wire(0) /=  '0') else type_cast_7788_wire_constant;
    -- logger for split-operator MUX_7799_inst flow-through 
    process(IMA88_7800) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_7799_inst:flowthrough inputs: " & " BITSEL_u8_u1_7794_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_7794_wire) & " type_cast_7796_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7796_wire_constant) & " type_cast_7798_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7798_wire_constant) & " outputs:" & " IMA88_7800= "  & Convert_SLV_To_Hex_String(IMA88_7800));
      --
    end process; 
    -- flow-through select operator MUX_7799_inst
    IMA88_7800 <= type_cast_7796_wire_constant when (BITSEL_u8_u1_7794_wire(0) /=  '0') else type_cast_7798_wire_constant;
    -- logger for split-operator MUX_7809_inst flow-through 
    process(IMA89_7810) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_7809_inst:flowthrough inputs: " & " BITSEL_u8_u1_7804_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_7804_wire) & " type_cast_7806_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7806_wire_constant) & " type_cast_7808_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7808_wire_constant) & " outputs:" & " IMA89_7810= "  & Convert_SLV_To_Hex_String(IMA89_7810));
      --
    end process; 
    -- flow-through select operator MUX_7809_inst
    IMA89_7810 <= type_cast_7806_wire_constant when (BITSEL_u8_u1_7804_wire(0) /=  '0') else type_cast_7808_wire_constant;
    -- logger for split-operator MUX_7819_inst flow-through 
    process(IMA90_7820) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_7819_inst:flowthrough inputs: " & " BITSEL_u8_u1_7814_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_7814_wire) & " type_cast_7816_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7816_wire_constant) & " type_cast_7818_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7818_wire_constant) & " outputs:" & " IMA90_7820= "  & Convert_SLV_To_Hex_String(IMA90_7820));
      --
    end process; 
    -- flow-through select operator MUX_7819_inst
    IMA90_7820 <= type_cast_7816_wire_constant when (BITSEL_u8_u1_7814_wire(0) /=  '0') else type_cast_7818_wire_constant;
    -- logger for split-operator MUX_7829_inst flow-through 
    process(IMA91_7830) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_7829_inst:flowthrough inputs: " & " BITSEL_u8_u1_7824_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_7824_wire) & " type_cast_7826_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7826_wire_constant) & " type_cast_7828_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7828_wire_constant) & " outputs:" & " IMA91_7830= "  & Convert_SLV_To_Hex_String(IMA91_7830));
      --
    end process; 
    -- flow-through select operator MUX_7829_inst
    IMA91_7830 <= type_cast_7826_wire_constant when (BITSEL_u8_u1_7824_wire(0) /=  '0') else type_cast_7828_wire_constant;
    -- logger for split-operator MUX_7839_inst flow-through 
    process(IMA92_7840) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_7839_inst:flowthrough inputs: " & " BITSEL_u8_u1_7834_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_7834_wire) & " type_cast_7836_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7836_wire_constant) & " type_cast_7838_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7838_wire_constant) & " outputs:" & " IMA92_7840= "  & Convert_SLV_To_Hex_String(IMA92_7840));
      --
    end process; 
    -- flow-through select operator MUX_7839_inst
    IMA92_7840 <= type_cast_7836_wire_constant when (BITSEL_u8_u1_7834_wire(0) /=  '0') else type_cast_7838_wire_constant;
    -- logger for split-operator MUX_7849_inst flow-through 
    process(IMA93_7850) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_7849_inst:flowthrough inputs: " & " BITSEL_u8_u1_7844_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_7844_wire) & " type_cast_7846_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7846_wire_constant) & " type_cast_7848_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7848_wire_constant) & " outputs:" & " IMA93_7850= "  & Convert_SLV_To_Hex_String(IMA93_7850));
      --
    end process; 
    -- flow-through select operator MUX_7849_inst
    IMA93_7850 <= type_cast_7846_wire_constant when (BITSEL_u8_u1_7844_wire(0) /=  '0') else type_cast_7848_wire_constant;
    -- logger for split-operator MUX_7859_inst flow-through 
    process(IMA94_7860) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_7859_inst:flowthrough inputs: " & " BITSEL_u8_u1_7854_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_7854_wire) & " type_cast_7856_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7856_wire_constant) & " type_cast_7858_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7858_wire_constant) & " outputs:" & " IMA94_7860= "  & Convert_SLV_To_Hex_String(IMA94_7860));
      --
    end process; 
    -- flow-through select operator MUX_7859_inst
    IMA94_7860 <= type_cast_7856_wire_constant when (BITSEL_u8_u1_7854_wire(0) /=  '0') else type_cast_7858_wire_constant;
    -- logger for split-operator MUX_7869_inst flow-through 
    process(IMA95_7870) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_7869_inst:flowthrough inputs: " & " BITSEL_u8_u1_7864_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_7864_wire) & " type_cast_7866_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7866_wire_constant) & " type_cast_7868_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7868_wire_constant) & " outputs:" & " IMA95_7870= "  & Convert_SLV_To_Hex_String(IMA95_7870));
      --
    end process; 
    -- flow-through select operator MUX_7869_inst
    IMA95_7870 <= type_cast_7866_wire_constant when (BITSEL_u8_u1_7864_wire(0) /=  '0') else type_cast_7868_wire_constant;
    -- logger for split-operator MUX_7879_inst flow-through 
    process(IMA96_7880) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_7879_inst:flowthrough inputs: " & " BITSEL_u8_u1_7874_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_7874_wire) & " type_cast_7876_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7876_wire_constant) & " type_cast_7878_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7878_wire_constant) & " outputs:" & " IMA96_7880= "  & Convert_SLV_To_Hex_String(IMA96_7880));
      --
    end process; 
    -- flow-through select operator MUX_7879_inst
    IMA96_7880 <= type_cast_7876_wire_constant when (BITSEL_u8_u1_7874_wire(0) /=  '0') else type_cast_7878_wire_constant;
    -- logger for split-operator MUX_7889_inst flow-through 
    process(IMA97_7890) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_7889_inst:flowthrough inputs: " & " BITSEL_u8_u1_7884_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_7884_wire) & " type_cast_7886_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7886_wire_constant) & " type_cast_7888_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7888_wire_constant) & " outputs:" & " IMA97_7890= "  & Convert_SLV_To_Hex_String(IMA97_7890));
      --
    end process; 
    -- flow-through select operator MUX_7889_inst
    IMA97_7890 <= type_cast_7886_wire_constant when (BITSEL_u8_u1_7884_wire(0) /=  '0') else type_cast_7888_wire_constant;
    -- logger for split-operator MUX_7899_inst flow-through 
    process(IMA98_7900) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_7899_inst:flowthrough inputs: " & " BITSEL_u8_u1_7894_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_7894_wire) & " type_cast_7896_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7896_wire_constant) & " type_cast_7898_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7898_wire_constant) & " outputs:" & " IMA98_7900= "  & Convert_SLV_To_Hex_String(IMA98_7900));
      --
    end process; 
    -- flow-through select operator MUX_7899_inst
    IMA98_7900 <= type_cast_7896_wire_constant when (BITSEL_u8_u1_7894_wire(0) /=  '0') else type_cast_7898_wire_constant;
    -- logger for split-operator MUX_7909_inst flow-through 
    process(IMA99_7910) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_7909_inst:flowthrough inputs: " & " BITSEL_u8_u1_7904_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_7904_wire) & " type_cast_7906_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7906_wire_constant) & " type_cast_7908_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7908_wire_constant) & " outputs:" & " IMA99_7910= "  & Convert_SLV_To_Hex_String(IMA99_7910));
      --
    end process; 
    -- flow-through select operator MUX_7909_inst
    IMA99_7910 <= type_cast_7906_wire_constant when (BITSEL_u8_u1_7904_wire(0) /=  '0') else type_cast_7908_wire_constant;
    -- logger for split-operator MUX_7919_inst flow-through 
    process(IMA100_7920) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_7919_inst:flowthrough inputs: " & " BITSEL_u8_u1_7914_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_7914_wire) & " type_cast_7916_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7916_wire_constant) & " type_cast_7918_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7918_wire_constant) & " outputs:" & " IMA100_7920= "  & Convert_SLV_To_Hex_String(IMA100_7920));
      --
    end process; 
    -- flow-through select operator MUX_7919_inst
    IMA100_7920 <= type_cast_7916_wire_constant when (BITSEL_u8_u1_7914_wire(0) /=  '0') else type_cast_7918_wire_constant;
    -- logger for split-operator MUX_7929_inst flow-through 
    process(IMA101_7930) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_7929_inst:flowthrough inputs: " & " BITSEL_u8_u1_7924_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_7924_wire) & " type_cast_7926_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7926_wire_constant) & " type_cast_7928_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7928_wire_constant) & " outputs:" & " IMA101_7930= "  & Convert_SLV_To_Hex_String(IMA101_7930));
      --
    end process; 
    -- flow-through select operator MUX_7929_inst
    IMA101_7930 <= type_cast_7926_wire_constant when (BITSEL_u8_u1_7924_wire(0) /=  '0') else type_cast_7928_wire_constant;
    -- logger for split-operator MUX_7939_inst flow-through 
    process(IMA102_7940) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_7939_inst:flowthrough inputs: " & " BITSEL_u8_u1_7934_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_7934_wire) & " type_cast_7936_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7936_wire_constant) & " type_cast_7938_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7938_wire_constant) & " outputs:" & " IMA102_7940= "  & Convert_SLV_To_Hex_String(IMA102_7940));
      --
    end process; 
    -- flow-through select operator MUX_7939_inst
    IMA102_7940 <= type_cast_7936_wire_constant when (BITSEL_u8_u1_7934_wire(0) /=  '0') else type_cast_7938_wire_constant;
    -- logger for split-operator MUX_7949_inst flow-through 
    process(IMA103_7950) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_7949_inst:flowthrough inputs: " & " BITSEL_u8_u1_7944_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_7944_wire) & " type_cast_7946_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7946_wire_constant) & " type_cast_7948_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7948_wire_constant) & " outputs:" & " IMA103_7950= "  & Convert_SLV_To_Hex_String(IMA103_7950));
      --
    end process; 
    -- flow-through select operator MUX_7949_inst
    IMA103_7950 <= type_cast_7946_wire_constant when (BITSEL_u8_u1_7944_wire(0) /=  '0') else type_cast_7948_wire_constant;
    -- logger for split-operator MUX_7959_inst flow-through 
    process(IMA104_7960) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_7959_inst:flowthrough inputs: " & " BITSEL_u8_u1_7954_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_7954_wire) & " type_cast_7956_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7956_wire_constant) & " type_cast_7958_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7958_wire_constant) & " outputs:" & " IMA104_7960= "  & Convert_SLV_To_Hex_String(IMA104_7960));
      --
    end process; 
    -- flow-through select operator MUX_7959_inst
    IMA104_7960 <= type_cast_7956_wire_constant when (BITSEL_u8_u1_7954_wire(0) /=  '0') else type_cast_7958_wire_constant;
    -- logger for split-operator MUX_7969_inst flow-through 
    process(IMA105_7970) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_7969_inst:flowthrough inputs: " & " BITSEL_u8_u1_7964_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_7964_wire) & " type_cast_7966_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7966_wire_constant) & " type_cast_7968_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7968_wire_constant) & " outputs:" & " IMA105_7970= "  & Convert_SLV_To_Hex_String(IMA105_7970));
      --
    end process; 
    -- flow-through select operator MUX_7969_inst
    IMA105_7970 <= type_cast_7966_wire_constant when (BITSEL_u8_u1_7964_wire(0) /=  '0') else type_cast_7968_wire_constant;
    -- logger for split-operator MUX_7979_inst flow-through 
    process(IMA106_7980) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_7979_inst:flowthrough inputs: " & " BITSEL_u8_u1_7974_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_7974_wire) & " type_cast_7976_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7976_wire_constant) & " type_cast_7978_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7978_wire_constant) & " outputs:" & " IMA106_7980= "  & Convert_SLV_To_Hex_String(IMA106_7980));
      --
    end process; 
    -- flow-through select operator MUX_7979_inst
    IMA106_7980 <= type_cast_7976_wire_constant when (BITSEL_u8_u1_7974_wire(0) /=  '0') else type_cast_7978_wire_constant;
    -- logger for split-operator MUX_7989_inst flow-through 
    process(IMA107_7990) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_7989_inst:flowthrough inputs: " & " BITSEL_u8_u1_7984_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_7984_wire) & " type_cast_7986_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7986_wire_constant) & " type_cast_7988_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7988_wire_constant) & " outputs:" & " IMA107_7990= "  & Convert_SLV_To_Hex_String(IMA107_7990));
      --
    end process; 
    -- flow-through select operator MUX_7989_inst
    IMA107_7990 <= type_cast_7986_wire_constant when (BITSEL_u8_u1_7984_wire(0) /=  '0') else type_cast_7988_wire_constant;
    -- logger for split-operator MUX_7999_inst flow-through 
    process(IMA108_8000) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_7999_inst:flowthrough inputs: " & " BITSEL_u8_u1_7994_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_7994_wire) & " type_cast_7996_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7996_wire_constant) & " type_cast_7998_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_7998_wire_constant) & " outputs:" & " IMA108_8000= "  & Convert_SLV_To_Hex_String(IMA108_8000));
      --
    end process; 
    -- flow-through select operator MUX_7999_inst
    IMA108_8000 <= type_cast_7996_wire_constant when (BITSEL_u8_u1_7994_wire(0) /=  '0') else type_cast_7998_wire_constant;
    -- logger for split-operator MUX_8009_inst flow-through 
    process(IMA109_8010) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8009_inst:flowthrough inputs: " & " BITSEL_u8_u1_8004_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8004_wire) & " type_cast_8006_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_8006_wire_constant) & " type_cast_8008_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_8008_wire_constant) & " outputs:" & " IMA109_8010= "  & Convert_SLV_To_Hex_String(IMA109_8010));
      --
    end process; 
    -- flow-through select operator MUX_8009_inst
    IMA109_8010 <= type_cast_8006_wire_constant when (BITSEL_u8_u1_8004_wire(0) /=  '0') else type_cast_8008_wire_constant;
    -- logger for split-operator MUX_8019_inst flow-through 
    process(IMA110_8020) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8019_inst:flowthrough inputs: " & " BITSEL_u8_u1_8014_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8014_wire) & " type_cast_8016_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_8016_wire_constant) & " type_cast_8018_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_8018_wire_constant) & " outputs:" & " IMA110_8020= "  & Convert_SLV_To_Hex_String(IMA110_8020));
      --
    end process; 
    -- flow-through select operator MUX_8019_inst
    IMA110_8020 <= type_cast_8016_wire_constant when (BITSEL_u8_u1_8014_wire(0) /=  '0') else type_cast_8018_wire_constant;
    -- logger for split-operator MUX_8029_inst flow-through 
    process(IMA111_8030) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8029_inst:flowthrough inputs: " & " BITSEL_u8_u1_8024_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8024_wire) & " type_cast_8026_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_8026_wire_constant) & " type_cast_8028_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_8028_wire_constant) & " outputs:" & " IMA111_8030= "  & Convert_SLV_To_Hex_String(IMA111_8030));
      --
    end process; 
    -- flow-through select operator MUX_8029_inst
    IMA111_8030 <= type_cast_8026_wire_constant when (BITSEL_u8_u1_8024_wire(0) /=  '0') else type_cast_8028_wire_constant;
    -- logger for split-operator MUX_8039_inst flow-through 
    process(IMA112_8040) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8039_inst:flowthrough inputs: " & " BITSEL_u8_u1_8034_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8034_wire) & " type_cast_8036_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_8036_wire_constant) & " type_cast_8038_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_8038_wire_constant) & " outputs:" & " IMA112_8040= "  & Convert_SLV_To_Hex_String(IMA112_8040));
      --
    end process; 
    -- flow-through select operator MUX_8039_inst
    IMA112_8040 <= type_cast_8036_wire_constant when (BITSEL_u8_u1_8034_wire(0) /=  '0') else type_cast_8038_wire_constant;
    -- logger for split-operator MUX_8049_inst flow-through 
    process(IMA113_8050) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8049_inst:flowthrough inputs: " & " BITSEL_u8_u1_8044_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8044_wire) & " type_cast_8046_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_8046_wire_constant) & " type_cast_8048_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_8048_wire_constant) & " outputs:" & " IMA113_8050= "  & Convert_SLV_To_Hex_String(IMA113_8050));
      --
    end process; 
    -- flow-through select operator MUX_8049_inst
    IMA113_8050 <= type_cast_8046_wire_constant when (BITSEL_u8_u1_8044_wire(0) /=  '0') else type_cast_8048_wire_constant;
    -- logger for split-operator MUX_8059_inst flow-through 
    process(IMA114_8060) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8059_inst:flowthrough inputs: " & " BITSEL_u8_u1_8054_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8054_wire) & " type_cast_8056_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_8056_wire_constant) & " type_cast_8058_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_8058_wire_constant) & " outputs:" & " IMA114_8060= "  & Convert_SLV_To_Hex_String(IMA114_8060));
      --
    end process; 
    -- flow-through select operator MUX_8059_inst
    IMA114_8060 <= type_cast_8056_wire_constant when (BITSEL_u8_u1_8054_wire(0) /=  '0') else type_cast_8058_wire_constant;
    -- logger for split-operator MUX_8069_inst flow-through 
    process(IMA115_8070) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8069_inst:flowthrough inputs: " & " BITSEL_u8_u1_8064_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8064_wire) & " type_cast_8066_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_8066_wire_constant) & " type_cast_8068_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_8068_wire_constant) & " outputs:" & " IMA115_8070= "  & Convert_SLV_To_Hex_String(IMA115_8070));
      --
    end process; 
    -- flow-through select operator MUX_8069_inst
    IMA115_8070 <= type_cast_8066_wire_constant when (BITSEL_u8_u1_8064_wire(0) /=  '0') else type_cast_8068_wire_constant;
    -- logger for split-operator MUX_8079_inst flow-through 
    process(IMA116_8080) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8079_inst:flowthrough inputs: " & " BITSEL_u8_u1_8074_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8074_wire) & " type_cast_8076_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_8076_wire_constant) & " type_cast_8078_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_8078_wire_constant) & " outputs:" & " IMA116_8080= "  & Convert_SLV_To_Hex_String(IMA116_8080));
      --
    end process; 
    -- flow-through select operator MUX_8079_inst
    IMA116_8080 <= type_cast_8076_wire_constant when (BITSEL_u8_u1_8074_wire(0) /=  '0') else type_cast_8078_wire_constant;
    -- logger for split-operator MUX_8089_inst flow-through 
    process(IMA117_8090) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8089_inst:flowthrough inputs: " & " BITSEL_u8_u1_8084_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8084_wire) & " type_cast_8086_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_8086_wire_constant) & " type_cast_8088_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_8088_wire_constant) & " outputs:" & " IMA117_8090= "  & Convert_SLV_To_Hex_String(IMA117_8090));
      --
    end process; 
    -- flow-through select operator MUX_8089_inst
    IMA117_8090 <= type_cast_8086_wire_constant when (BITSEL_u8_u1_8084_wire(0) /=  '0') else type_cast_8088_wire_constant;
    -- logger for split-operator MUX_8099_inst flow-through 
    process(IMA118_8100) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8099_inst:flowthrough inputs: " & " BITSEL_u8_u1_8094_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8094_wire) & " type_cast_8096_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_8096_wire_constant) & " type_cast_8098_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_8098_wire_constant) & " outputs:" & " IMA118_8100= "  & Convert_SLV_To_Hex_String(IMA118_8100));
      --
    end process; 
    -- flow-through select operator MUX_8099_inst
    IMA118_8100 <= type_cast_8096_wire_constant when (BITSEL_u8_u1_8094_wire(0) /=  '0') else type_cast_8098_wire_constant;
    -- logger for split-operator MUX_8109_inst flow-through 
    process(IMA119_8110) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8109_inst:flowthrough inputs: " & " BITSEL_u8_u1_8104_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8104_wire) & " type_cast_8106_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_8106_wire_constant) & " type_cast_8108_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_8108_wire_constant) & " outputs:" & " IMA119_8110= "  & Convert_SLV_To_Hex_String(IMA119_8110));
      --
    end process; 
    -- flow-through select operator MUX_8109_inst
    IMA119_8110 <= type_cast_8106_wire_constant when (BITSEL_u8_u1_8104_wire(0) /=  '0') else type_cast_8108_wire_constant;
    -- logger for split-operator MUX_8119_inst flow-through 
    process(IMA120_8120) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8119_inst:flowthrough inputs: " & " BITSEL_u8_u1_8114_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8114_wire) & " type_cast_8116_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_8116_wire_constant) & " type_cast_8118_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_8118_wire_constant) & " outputs:" & " IMA120_8120= "  & Convert_SLV_To_Hex_String(IMA120_8120));
      --
    end process; 
    -- flow-through select operator MUX_8119_inst
    IMA120_8120 <= type_cast_8116_wire_constant when (BITSEL_u8_u1_8114_wire(0) /=  '0') else type_cast_8118_wire_constant;
    -- logger for split-operator MUX_8129_inst flow-through 
    process(IMA121_8130) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8129_inst:flowthrough inputs: " & " BITSEL_u8_u1_8124_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8124_wire) & " type_cast_8126_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_8126_wire_constant) & " type_cast_8128_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_8128_wire_constant) & " outputs:" & " IMA121_8130= "  & Convert_SLV_To_Hex_String(IMA121_8130));
      --
    end process; 
    -- flow-through select operator MUX_8129_inst
    IMA121_8130 <= type_cast_8126_wire_constant when (BITSEL_u8_u1_8124_wire(0) /=  '0') else type_cast_8128_wire_constant;
    -- logger for split-operator MUX_8139_inst flow-through 
    process(IMA122_8140) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8139_inst:flowthrough inputs: " & " BITSEL_u8_u1_8134_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8134_wire) & " type_cast_8136_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_8136_wire_constant) & " type_cast_8138_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_8138_wire_constant) & " outputs:" & " IMA122_8140= "  & Convert_SLV_To_Hex_String(IMA122_8140));
      --
    end process; 
    -- flow-through select operator MUX_8139_inst
    IMA122_8140 <= type_cast_8136_wire_constant when (BITSEL_u8_u1_8134_wire(0) /=  '0') else type_cast_8138_wire_constant;
    -- logger for split-operator MUX_8149_inst flow-through 
    process(IMA123_8150) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8149_inst:flowthrough inputs: " & " BITSEL_u8_u1_8144_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8144_wire) & " type_cast_8146_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_8146_wire_constant) & " type_cast_8148_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_8148_wire_constant) & " outputs:" & " IMA123_8150= "  & Convert_SLV_To_Hex_String(IMA123_8150));
      --
    end process; 
    -- flow-through select operator MUX_8149_inst
    IMA123_8150 <= type_cast_8146_wire_constant when (BITSEL_u8_u1_8144_wire(0) /=  '0') else type_cast_8148_wire_constant;
    -- logger for split-operator MUX_8159_inst flow-through 
    process(IMA124_8160) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8159_inst:flowthrough inputs: " & " BITSEL_u8_u1_8154_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8154_wire) & " type_cast_8156_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_8156_wire_constant) & " type_cast_8158_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_8158_wire_constant) & " outputs:" & " IMA124_8160= "  & Convert_SLV_To_Hex_String(IMA124_8160));
      --
    end process; 
    -- flow-through select operator MUX_8159_inst
    IMA124_8160 <= type_cast_8156_wire_constant when (BITSEL_u8_u1_8154_wire(0) /=  '0') else type_cast_8158_wire_constant;
    -- logger for split-operator MUX_8169_inst flow-through 
    process(IMA125_8170) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8169_inst:flowthrough inputs: " & " BITSEL_u8_u1_8164_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8164_wire) & " type_cast_8166_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_8166_wire_constant) & " type_cast_8168_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_8168_wire_constant) & " outputs:" & " IMA125_8170= "  & Convert_SLV_To_Hex_String(IMA125_8170));
      --
    end process; 
    -- flow-through select operator MUX_8169_inst
    IMA125_8170 <= type_cast_8166_wire_constant when (BITSEL_u8_u1_8164_wire(0) /=  '0') else type_cast_8168_wire_constant;
    -- logger for split-operator MUX_8179_inst flow-through 
    process(IMA126_8180) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8179_inst:flowthrough inputs: " & " BITSEL_u8_u1_8174_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8174_wire) & " type_cast_8176_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_8176_wire_constant) & " type_cast_8178_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_8178_wire_constant) & " outputs:" & " IMA126_8180= "  & Convert_SLV_To_Hex_String(IMA126_8180));
      --
    end process; 
    -- flow-through select operator MUX_8179_inst
    IMA126_8180 <= type_cast_8176_wire_constant when (BITSEL_u8_u1_8174_wire(0) /=  '0') else type_cast_8178_wire_constant;
    -- logger for split-operator MUX_8189_inst flow-through 
    process(IMA127_8190) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8189_inst:flowthrough inputs: " & " BITSEL_u8_u1_8184_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8184_wire) & " type_cast_8186_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_8186_wire_constant) & " type_cast_8188_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_8188_wire_constant) & " outputs:" & " IMA127_8190= "  & Convert_SLV_To_Hex_String(IMA127_8190));
      --
    end process; 
    -- flow-through select operator MUX_8189_inst
    IMA127_8190 <= type_cast_8186_wire_constant when (BITSEL_u8_u1_8184_wire(0) /=  '0') else type_cast_8188_wire_constant;
    -- logger for split-operator MUX_8197_inst flow-through 
    process(IMB0_8198) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8197_inst:flowthrough inputs: " & " BITSEL_u8_u1_8194_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8194_wire) & " IMA1_6930 = "& Convert_SLV_To_Hex_String(IMA1_6930) & " IMA0_6920 = "& Convert_SLV_To_Hex_String(IMA0_6920) & " outputs:" & " IMB0_8198= "  & Convert_SLV_To_Hex_String(IMB0_8198));
      --
    end process; 
    -- flow-through select operator MUX_8197_inst
    IMB0_8198 <= IMA1_6930 when (BITSEL_u8_u1_8194_wire(0) /=  '0') else IMA0_6920;
    -- logger for split-operator MUX_8205_inst flow-through 
    process(IMB1_8206) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8205_inst:flowthrough inputs: " & " BITSEL_u8_u1_8202_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8202_wire) & " IMA3_6950 = "& Convert_SLV_To_Hex_String(IMA3_6950) & " IMA2_6940 = "& Convert_SLV_To_Hex_String(IMA2_6940) & " outputs:" & " IMB1_8206= "  & Convert_SLV_To_Hex_String(IMB1_8206));
      --
    end process; 
    -- flow-through select operator MUX_8205_inst
    IMB1_8206 <= IMA3_6950 when (BITSEL_u8_u1_8202_wire(0) /=  '0') else IMA2_6940;
    -- logger for split-operator MUX_8213_inst flow-through 
    process(IMB2_8214) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8213_inst:flowthrough inputs: " & " BITSEL_u8_u1_8210_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8210_wire) & " IMA5_6970 = "& Convert_SLV_To_Hex_String(IMA5_6970) & " IMA4_6960 = "& Convert_SLV_To_Hex_String(IMA4_6960) & " outputs:" & " IMB2_8214= "  & Convert_SLV_To_Hex_String(IMB2_8214));
      --
    end process; 
    -- flow-through select operator MUX_8213_inst
    IMB2_8214 <= IMA5_6970 when (BITSEL_u8_u1_8210_wire(0) /=  '0') else IMA4_6960;
    -- logger for split-operator MUX_8221_inst flow-through 
    process(IMB3_8222) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8221_inst:flowthrough inputs: " & " BITSEL_u8_u1_8218_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8218_wire) & " IMA7_6990 = "& Convert_SLV_To_Hex_String(IMA7_6990) & " IMA6_6980 = "& Convert_SLV_To_Hex_String(IMA6_6980) & " outputs:" & " IMB3_8222= "  & Convert_SLV_To_Hex_String(IMB3_8222));
      --
    end process; 
    -- flow-through select operator MUX_8221_inst
    IMB3_8222 <= IMA7_6990 when (BITSEL_u8_u1_8218_wire(0) /=  '0') else IMA6_6980;
    -- logger for split-operator MUX_8229_inst flow-through 
    process(IMB4_8230) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8229_inst:flowthrough inputs: " & " BITSEL_u8_u1_8226_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8226_wire) & " IMA9_7010 = "& Convert_SLV_To_Hex_String(IMA9_7010) & " IMA8_7000 = "& Convert_SLV_To_Hex_String(IMA8_7000) & " outputs:" & " IMB4_8230= "  & Convert_SLV_To_Hex_String(IMB4_8230));
      --
    end process; 
    -- flow-through select operator MUX_8229_inst
    IMB4_8230 <= IMA9_7010 when (BITSEL_u8_u1_8226_wire(0) /=  '0') else IMA8_7000;
    -- logger for split-operator MUX_8237_inst flow-through 
    process(IMB5_8238) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8237_inst:flowthrough inputs: " & " BITSEL_u8_u1_8234_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8234_wire) & " IMA11_7030 = "& Convert_SLV_To_Hex_String(IMA11_7030) & " IMA10_7020 = "& Convert_SLV_To_Hex_String(IMA10_7020) & " outputs:" & " IMB5_8238= "  & Convert_SLV_To_Hex_String(IMB5_8238));
      --
    end process; 
    -- flow-through select operator MUX_8237_inst
    IMB5_8238 <= IMA11_7030 when (BITSEL_u8_u1_8234_wire(0) /=  '0') else IMA10_7020;
    -- logger for split-operator MUX_8245_inst flow-through 
    process(IMB6_8246) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8245_inst:flowthrough inputs: " & " BITSEL_u8_u1_8242_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8242_wire) & " IMA13_7050 = "& Convert_SLV_To_Hex_String(IMA13_7050) & " IMA12_7040 = "& Convert_SLV_To_Hex_String(IMA12_7040) & " outputs:" & " IMB6_8246= "  & Convert_SLV_To_Hex_String(IMB6_8246));
      --
    end process; 
    -- flow-through select operator MUX_8245_inst
    IMB6_8246 <= IMA13_7050 when (BITSEL_u8_u1_8242_wire(0) /=  '0') else IMA12_7040;
    -- logger for split-operator MUX_8253_inst flow-through 
    process(IMB7_8254) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8253_inst:flowthrough inputs: " & " BITSEL_u8_u1_8250_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8250_wire) & " IMA15_7070 = "& Convert_SLV_To_Hex_String(IMA15_7070) & " IMA14_7060 = "& Convert_SLV_To_Hex_String(IMA14_7060) & " outputs:" & " IMB7_8254= "  & Convert_SLV_To_Hex_String(IMB7_8254));
      --
    end process; 
    -- flow-through select operator MUX_8253_inst
    IMB7_8254 <= IMA15_7070 when (BITSEL_u8_u1_8250_wire(0) /=  '0') else IMA14_7060;
    -- logger for split-operator MUX_8261_inst flow-through 
    process(IMB8_8262) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8261_inst:flowthrough inputs: " & " BITSEL_u8_u1_8258_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8258_wire) & " IMA17_7090 = "& Convert_SLV_To_Hex_String(IMA17_7090) & " IMA16_7080 = "& Convert_SLV_To_Hex_String(IMA16_7080) & " outputs:" & " IMB8_8262= "  & Convert_SLV_To_Hex_String(IMB8_8262));
      --
    end process; 
    -- flow-through select operator MUX_8261_inst
    IMB8_8262 <= IMA17_7090 when (BITSEL_u8_u1_8258_wire(0) /=  '0') else IMA16_7080;
    -- logger for split-operator MUX_8269_inst flow-through 
    process(IMB9_8270) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8269_inst:flowthrough inputs: " & " BITSEL_u8_u1_8266_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8266_wire) & " IMA19_7110 = "& Convert_SLV_To_Hex_String(IMA19_7110) & " IMA18_7100 = "& Convert_SLV_To_Hex_String(IMA18_7100) & " outputs:" & " IMB9_8270= "  & Convert_SLV_To_Hex_String(IMB9_8270));
      --
    end process; 
    -- flow-through select operator MUX_8269_inst
    IMB9_8270 <= IMA19_7110 when (BITSEL_u8_u1_8266_wire(0) /=  '0') else IMA18_7100;
    -- logger for split-operator MUX_8277_inst flow-through 
    process(IMB10_8278) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8277_inst:flowthrough inputs: " & " BITSEL_u8_u1_8274_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8274_wire) & " IMA21_7130 = "& Convert_SLV_To_Hex_String(IMA21_7130) & " IMA20_7120 = "& Convert_SLV_To_Hex_String(IMA20_7120) & " outputs:" & " IMB10_8278= "  & Convert_SLV_To_Hex_String(IMB10_8278));
      --
    end process; 
    -- flow-through select operator MUX_8277_inst
    IMB10_8278 <= IMA21_7130 when (BITSEL_u8_u1_8274_wire(0) /=  '0') else IMA20_7120;
    -- logger for split-operator MUX_8285_inst flow-through 
    process(IMB11_8286) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8285_inst:flowthrough inputs: " & " BITSEL_u8_u1_8282_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8282_wire) & " IMA23_7150 = "& Convert_SLV_To_Hex_String(IMA23_7150) & " IMA22_7140 = "& Convert_SLV_To_Hex_String(IMA22_7140) & " outputs:" & " IMB11_8286= "  & Convert_SLV_To_Hex_String(IMB11_8286));
      --
    end process; 
    -- flow-through select operator MUX_8285_inst
    IMB11_8286 <= IMA23_7150 when (BITSEL_u8_u1_8282_wire(0) /=  '0') else IMA22_7140;
    -- logger for split-operator MUX_8293_inst flow-through 
    process(IMB12_8294) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8293_inst:flowthrough inputs: " & " BITSEL_u8_u1_8290_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8290_wire) & " IMA25_7170 = "& Convert_SLV_To_Hex_String(IMA25_7170) & " IMA24_7160 = "& Convert_SLV_To_Hex_String(IMA24_7160) & " outputs:" & " IMB12_8294= "  & Convert_SLV_To_Hex_String(IMB12_8294));
      --
    end process; 
    -- flow-through select operator MUX_8293_inst
    IMB12_8294 <= IMA25_7170 when (BITSEL_u8_u1_8290_wire(0) /=  '0') else IMA24_7160;
    -- logger for split-operator MUX_8301_inst flow-through 
    process(IMB13_8302) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8301_inst:flowthrough inputs: " & " BITSEL_u8_u1_8298_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8298_wire) & " IMA27_7190 = "& Convert_SLV_To_Hex_String(IMA27_7190) & " IMA26_7180 = "& Convert_SLV_To_Hex_String(IMA26_7180) & " outputs:" & " IMB13_8302= "  & Convert_SLV_To_Hex_String(IMB13_8302));
      --
    end process; 
    -- flow-through select operator MUX_8301_inst
    IMB13_8302 <= IMA27_7190 when (BITSEL_u8_u1_8298_wire(0) /=  '0') else IMA26_7180;
    -- logger for split-operator MUX_8309_inst flow-through 
    process(IMB14_8310) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8309_inst:flowthrough inputs: " & " BITSEL_u8_u1_8306_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8306_wire) & " IMA29_7210 = "& Convert_SLV_To_Hex_String(IMA29_7210) & " IMA28_7200 = "& Convert_SLV_To_Hex_String(IMA28_7200) & " outputs:" & " IMB14_8310= "  & Convert_SLV_To_Hex_String(IMB14_8310));
      --
    end process; 
    -- flow-through select operator MUX_8309_inst
    IMB14_8310 <= IMA29_7210 when (BITSEL_u8_u1_8306_wire(0) /=  '0') else IMA28_7200;
    -- logger for split-operator MUX_8317_inst flow-through 
    process(IMB15_8318) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8317_inst:flowthrough inputs: " & " BITSEL_u8_u1_8314_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8314_wire) & " IMA31_7230 = "& Convert_SLV_To_Hex_String(IMA31_7230) & " IMA30_7220 = "& Convert_SLV_To_Hex_String(IMA30_7220) & " outputs:" & " IMB15_8318= "  & Convert_SLV_To_Hex_String(IMB15_8318));
      --
    end process; 
    -- flow-through select operator MUX_8317_inst
    IMB15_8318 <= IMA31_7230 when (BITSEL_u8_u1_8314_wire(0) /=  '0') else IMA30_7220;
    -- logger for split-operator MUX_8325_inst flow-through 
    process(IMB16_8326) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8325_inst:flowthrough inputs: " & " BITSEL_u8_u1_8322_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8322_wire) & " IMA33_7250 = "& Convert_SLV_To_Hex_String(IMA33_7250) & " IMA32_7240 = "& Convert_SLV_To_Hex_String(IMA32_7240) & " outputs:" & " IMB16_8326= "  & Convert_SLV_To_Hex_String(IMB16_8326));
      --
    end process; 
    -- flow-through select operator MUX_8325_inst
    IMB16_8326 <= IMA33_7250 when (BITSEL_u8_u1_8322_wire(0) /=  '0') else IMA32_7240;
    -- logger for split-operator MUX_8333_inst flow-through 
    process(IMB17_8334) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8333_inst:flowthrough inputs: " & " BITSEL_u8_u1_8330_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8330_wire) & " IMA35_7270 = "& Convert_SLV_To_Hex_String(IMA35_7270) & " IMA34_7260 = "& Convert_SLV_To_Hex_String(IMA34_7260) & " outputs:" & " IMB17_8334= "  & Convert_SLV_To_Hex_String(IMB17_8334));
      --
    end process; 
    -- flow-through select operator MUX_8333_inst
    IMB17_8334 <= IMA35_7270 when (BITSEL_u8_u1_8330_wire(0) /=  '0') else IMA34_7260;
    -- logger for split-operator MUX_8341_inst flow-through 
    process(IMB18_8342) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8341_inst:flowthrough inputs: " & " BITSEL_u8_u1_8338_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8338_wire) & " IMA37_7290 = "& Convert_SLV_To_Hex_String(IMA37_7290) & " IMA36_7280 = "& Convert_SLV_To_Hex_String(IMA36_7280) & " outputs:" & " IMB18_8342= "  & Convert_SLV_To_Hex_String(IMB18_8342));
      --
    end process; 
    -- flow-through select operator MUX_8341_inst
    IMB18_8342 <= IMA37_7290 when (BITSEL_u8_u1_8338_wire(0) /=  '0') else IMA36_7280;
    -- logger for split-operator MUX_8349_inst flow-through 
    process(IMB19_8350) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8349_inst:flowthrough inputs: " & " BITSEL_u8_u1_8346_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8346_wire) & " IMA39_7310 = "& Convert_SLV_To_Hex_String(IMA39_7310) & " IMA38_7300 = "& Convert_SLV_To_Hex_String(IMA38_7300) & " outputs:" & " IMB19_8350= "  & Convert_SLV_To_Hex_String(IMB19_8350));
      --
    end process; 
    -- flow-through select operator MUX_8349_inst
    IMB19_8350 <= IMA39_7310 when (BITSEL_u8_u1_8346_wire(0) /=  '0') else IMA38_7300;
    -- logger for split-operator MUX_8357_inst flow-through 
    process(IMB20_8358) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8357_inst:flowthrough inputs: " & " BITSEL_u8_u1_8354_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8354_wire) & " IMA41_7330 = "& Convert_SLV_To_Hex_String(IMA41_7330) & " IMA40_7320 = "& Convert_SLV_To_Hex_String(IMA40_7320) & " outputs:" & " IMB20_8358= "  & Convert_SLV_To_Hex_String(IMB20_8358));
      --
    end process; 
    -- flow-through select operator MUX_8357_inst
    IMB20_8358 <= IMA41_7330 when (BITSEL_u8_u1_8354_wire(0) /=  '0') else IMA40_7320;
    -- logger for split-operator MUX_8365_inst flow-through 
    process(IMB21_8366) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8365_inst:flowthrough inputs: " & " BITSEL_u8_u1_8362_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8362_wire) & " IMA43_7350 = "& Convert_SLV_To_Hex_String(IMA43_7350) & " IMA42_7340 = "& Convert_SLV_To_Hex_String(IMA42_7340) & " outputs:" & " IMB21_8366= "  & Convert_SLV_To_Hex_String(IMB21_8366));
      --
    end process; 
    -- flow-through select operator MUX_8365_inst
    IMB21_8366 <= IMA43_7350 when (BITSEL_u8_u1_8362_wire(0) /=  '0') else IMA42_7340;
    -- logger for split-operator MUX_8373_inst flow-through 
    process(IMB22_8374) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8373_inst:flowthrough inputs: " & " BITSEL_u8_u1_8370_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8370_wire) & " IMA45_7370 = "& Convert_SLV_To_Hex_String(IMA45_7370) & " IMA44_7360 = "& Convert_SLV_To_Hex_String(IMA44_7360) & " outputs:" & " IMB22_8374= "  & Convert_SLV_To_Hex_String(IMB22_8374));
      --
    end process; 
    -- flow-through select operator MUX_8373_inst
    IMB22_8374 <= IMA45_7370 when (BITSEL_u8_u1_8370_wire(0) /=  '0') else IMA44_7360;
    -- logger for split-operator MUX_8381_inst flow-through 
    process(IMB23_8382) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8381_inst:flowthrough inputs: " & " BITSEL_u8_u1_8378_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8378_wire) & " IMA47_7390 = "& Convert_SLV_To_Hex_String(IMA47_7390) & " IMA46_7380 = "& Convert_SLV_To_Hex_String(IMA46_7380) & " outputs:" & " IMB23_8382= "  & Convert_SLV_To_Hex_String(IMB23_8382));
      --
    end process; 
    -- flow-through select operator MUX_8381_inst
    IMB23_8382 <= IMA47_7390 when (BITSEL_u8_u1_8378_wire(0) /=  '0') else IMA46_7380;
    -- logger for split-operator MUX_8389_inst flow-through 
    process(IMB24_8390) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8389_inst:flowthrough inputs: " & " BITSEL_u8_u1_8386_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8386_wire) & " IMA49_7410 = "& Convert_SLV_To_Hex_String(IMA49_7410) & " IMA48_7400 = "& Convert_SLV_To_Hex_String(IMA48_7400) & " outputs:" & " IMB24_8390= "  & Convert_SLV_To_Hex_String(IMB24_8390));
      --
    end process; 
    -- flow-through select operator MUX_8389_inst
    IMB24_8390 <= IMA49_7410 when (BITSEL_u8_u1_8386_wire(0) /=  '0') else IMA48_7400;
    -- logger for split-operator MUX_8397_inst flow-through 
    process(IMB25_8398) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8397_inst:flowthrough inputs: " & " BITSEL_u8_u1_8394_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8394_wire) & " IMA51_7430 = "& Convert_SLV_To_Hex_String(IMA51_7430) & " IMA50_7420 = "& Convert_SLV_To_Hex_String(IMA50_7420) & " outputs:" & " IMB25_8398= "  & Convert_SLV_To_Hex_String(IMB25_8398));
      --
    end process; 
    -- flow-through select operator MUX_8397_inst
    IMB25_8398 <= IMA51_7430 when (BITSEL_u8_u1_8394_wire(0) /=  '0') else IMA50_7420;
    -- logger for split-operator MUX_8405_inst flow-through 
    process(IMB26_8406) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8405_inst:flowthrough inputs: " & " BITSEL_u8_u1_8402_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8402_wire) & " IMA53_7450 = "& Convert_SLV_To_Hex_String(IMA53_7450) & " IMA52_7440 = "& Convert_SLV_To_Hex_String(IMA52_7440) & " outputs:" & " IMB26_8406= "  & Convert_SLV_To_Hex_String(IMB26_8406));
      --
    end process; 
    -- flow-through select operator MUX_8405_inst
    IMB26_8406 <= IMA53_7450 when (BITSEL_u8_u1_8402_wire(0) /=  '0') else IMA52_7440;
    -- logger for split-operator MUX_8413_inst flow-through 
    process(IMB27_8414) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8413_inst:flowthrough inputs: " & " BITSEL_u8_u1_8410_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8410_wire) & " IMA55_7470 = "& Convert_SLV_To_Hex_String(IMA55_7470) & " IMA54_7460 = "& Convert_SLV_To_Hex_String(IMA54_7460) & " outputs:" & " IMB27_8414= "  & Convert_SLV_To_Hex_String(IMB27_8414));
      --
    end process; 
    -- flow-through select operator MUX_8413_inst
    IMB27_8414 <= IMA55_7470 when (BITSEL_u8_u1_8410_wire(0) /=  '0') else IMA54_7460;
    -- logger for split-operator MUX_8421_inst flow-through 
    process(IMB28_8422) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8421_inst:flowthrough inputs: " & " BITSEL_u8_u1_8418_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8418_wire) & " IMA57_7490 = "& Convert_SLV_To_Hex_String(IMA57_7490) & " IMA56_7480 = "& Convert_SLV_To_Hex_String(IMA56_7480) & " outputs:" & " IMB28_8422= "  & Convert_SLV_To_Hex_String(IMB28_8422));
      --
    end process; 
    -- flow-through select operator MUX_8421_inst
    IMB28_8422 <= IMA57_7490 when (BITSEL_u8_u1_8418_wire(0) /=  '0') else IMA56_7480;
    -- logger for split-operator MUX_8429_inst flow-through 
    process(IMB29_8430) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8429_inst:flowthrough inputs: " & " BITSEL_u8_u1_8426_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8426_wire) & " IMA59_7510 = "& Convert_SLV_To_Hex_String(IMA59_7510) & " IMA58_7500 = "& Convert_SLV_To_Hex_String(IMA58_7500) & " outputs:" & " IMB29_8430= "  & Convert_SLV_To_Hex_String(IMB29_8430));
      --
    end process; 
    -- flow-through select operator MUX_8429_inst
    IMB29_8430 <= IMA59_7510 when (BITSEL_u8_u1_8426_wire(0) /=  '0') else IMA58_7500;
    -- logger for split-operator MUX_8437_inst flow-through 
    process(IMB30_8438) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8437_inst:flowthrough inputs: " & " BITSEL_u8_u1_8434_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8434_wire) & " IMA61_7530 = "& Convert_SLV_To_Hex_String(IMA61_7530) & " IMA60_7520 = "& Convert_SLV_To_Hex_String(IMA60_7520) & " outputs:" & " IMB30_8438= "  & Convert_SLV_To_Hex_String(IMB30_8438));
      --
    end process; 
    -- flow-through select operator MUX_8437_inst
    IMB30_8438 <= IMA61_7530 when (BITSEL_u8_u1_8434_wire(0) /=  '0') else IMA60_7520;
    -- logger for split-operator MUX_8445_inst flow-through 
    process(IMB31_8446) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8445_inst:flowthrough inputs: " & " BITSEL_u8_u1_8442_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8442_wire) & " IMA63_7550 = "& Convert_SLV_To_Hex_String(IMA63_7550) & " IMA62_7540 = "& Convert_SLV_To_Hex_String(IMA62_7540) & " outputs:" & " IMB31_8446= "  & Convert_SLV_To_Hex_String(IMB31_8446));
      --
    end process; 
    -- flow-through select operator MUX_8445_inst
    IMB31_8446 <= IMA63_7550 when (BITSEL_u8_u1_8442_wire(0) /=  '0') else IMA62_7540;
    -- logger for split-operator MUX_8453_inst flow-through 
    process(IMB32_8454) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8453_inst:flowthrough inputs: " & " BITSEL_u8_u1_8450_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8450_wire) & " IMA65_7570 = "& Convert_SLV_To_Hex_String(IMA65_7570) & " IMA64_7560 = "& Convert_SLV_To_Hex_String(IMA64_7560) & " outputs:" & " IMB32_8454= "  & Convert_SLV_To_Hex_String(IMB32_8454));
      --
    end process; 
    -- flow-through select operator MUX_8453_inst
    IMB32_8454 <= IMA65_7570 when (BITSEL_u8_u1_8450_wire(0) /=  '0') else IMA64_7560;
    -- logger for split-operator MUX_8461_inst flow-through 
    process(IMB33_8462) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8461_inst:flowthrough inputs: " & " BITSEL_u8_u1_8458_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8458_wire) & " IMA67_7590 = "& Convert_SLV_To_Hex_String(IMA67_7590) & " IMA66_7580 = "& Convert_SLV_To_Hex_String(IMA66_7580) & " outputs:" & " IMB33_8462= "  & Convert_SLV_To_Hex_String(IMB33_8462));
      --
    end process; 
    -- flow-through select operator MUX_8461_inst
    IMB33_8462 <= IMA67_7590 when (BITSEL_u8_u1_8458_wire(0) /=  '0') else IMA66_7580;
    -- logger for split-operator MUX_8469_inst flow-through 
    process(IMB34_8470) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8469_inst:flowthrough inputs: " & " BITSEL_u8_u1_8466_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8466_wire) & " IMA69_7610 = "& Convert_SLV_To_Hex_String(IMA69_7610) & " IMA68_7600 = "& Convert_SLV_To_Hex_String(IMA68_7600) & " outputs:" & " IMB34_8470= "  & Convert_SLV_To_Hex_String(IMB34_8470));
      --
    end process; 
    -- flow-through select operator MUX_8469_inst
    IMB34_8470 <= IMA69_7610 when (BITSEL_u8_u1_8466_wire(0) /=  '0') else IMA68_7600;
    -- logger for split-operator MUX_8477_inst flow-through 
    process(IMB35_8478) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8477_inst:flowthrough inputs: " & " BITSEL_u8_u1_8474_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8474_wire) & " IMA71_7630 = "& Convert_SLV_To_Hex_String(IMA71_7630) & " IMA70_7620 = "& Convert_SLV_To_Hex_String(IMA70_7620) & " outputs:" & " IMB35_8478= "  & Convert_SLV_To_Hex_String(IMB35_8478));
      --
    end process; 
    -- flow-through select operator MUX_8477_inst
    IMB35_8478 <= IMA71_7630 when (BITSEL_u8_u1_8474_wire(0) /=  '0') else IMA70_7620;
    -- logger for split-operator MUX_8485_inst flow-through 
    process(IMB36_8486) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8485_inst:flowthrough inputs: " & " BITSEL_u8_u1_8482_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8482_wire) & " IMA73_7650 = "& Convert_SLV_To_Hex_String(IMA73_7650) & " IMA72_7640 = "& Convert_SLV_To_Hex_String(IMA72_7640) & " outputs:" & " IMB36_8486= "  & Convert_SLV_To_Hex_String(IMB36_8486));
      --
    end process; 
    -- flow-through select operator MUX_8485_inst
    IMB36_8486 <= IMA73_7650 when (BITSEL_u8_u1_8482_wire(0) /=  '0') else IMA72_7640;
    -- logger for split-operator MUX_8493_inst flow-through 
    process(IMB37_8494) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8493_inst:flowthrough inputs: " & " BITSEL_u8_u1_8490_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8490_wire) & " IMA75_7670 = "& Convert_SLV_To_Hex_String(IMA75_7670) & " IMA74_7660 = "& Convert_SLV_To_Hex_String(IMA74_7660) & " outputs:" & " IMB37_8494= "  & Convert_SLV_To_Hex_String(IMB37_8494));
      --
    end process; 
    -- flow-through select operator MUX_8493_inst
    IMB37_8494 <= IMA75_7670 when (BITSEL_u8_u1_8490_wire(0) /=  '0') else IMA74_7660;
    -- logger for split-operator MUX_8501_inst flow-through 
    process(IMB38_8502) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8501_inst:flowthrough inputs: " & " BITSEL_u8_u1_8498_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8498_wire) & " IMA77_7690 = "& Convert_SLV_To_Hex_String(IMA77_7690) & " IMA76_7680 = "& Convert_SLV_To_Hex_String(IMA76_7680) & " outputs:" & " IMB38_8502= "  & Convert_SLV_To_Hex_String(IMB38_8502));
      --
    end process; 
    -- flow-through select operator MUX_8501_inst
    IMB38_8502 <= IMA77_7690 when (BITSEL_u8_u1_8498_wire(0) /=  '0') else IMA76_7680;
    -- logger for split-operator MUX_8509_inst flow-through 
    process(IMB39_8510) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8509_inst:flowthrough inputs: " & " BITSEL_u8_u1_8506_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8506_wire) & " IMA79_7710 = "& Convert_SLV_To_Hex_String(IMA79_7710) & " IMA78_7700 = "& Convert_SLV_To_Hex_String(IMA78_7700) & " outputs:" & " IMB39_8510= "  & Convert_SLV_To_Hex_String(IMB39_8510));
      --
    end process; 
    -- flow-through select operator MUX_8509_inst
    IMB39_8510 <= IMA79_7710 when (BITSEL_u8_u1_8506_wire(0) /=  '0') else IMA78_7700;
    -- logger for split-operator MUX_8517_inst flow-through 
    process(IMB40_8518) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8517_inst:flowthrough inputs: " & " BITSEL_u8_u1_8514_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8514_wire) & " IMA81_7730 = "& Convert_SLV_To_Hex_String(IMA81_7730) & " IMA80_7720 = "& Convert_SLV_To_Hex_String(IMA80_7720) & " outputs:" & " IMB40_8518= "  & Convert_SLV_To_Hex_String(IMB40_8518));
      --
    end process; 
    -- flow-through select operator MUX_8517_inst
    IMB40_8518 <= IMA81_7730 when (BITSEL_u8_u1_8514_wire(0) /=  '0') else IMA80_7720;
    -- logger for split-operator MUX_8525_inst flow-through 
    process(IMB41_8526) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8525_inst:flowthrough inputs: " & " BITSEL_u8_u1_8522_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8522_wire) & " IMA83_7750 = "& Convert_SLV_To_Hex_String(IMA83_7750) & " IMA82_7740 = "& Convert_SLV_To_Hex_String(IMA82_7740) & " outputs:" & " IMB41_8526= "  & Convert_SLV_To_Hex_String(IMB41_8526));
      --
    end process; 
    -- flow-through select operator MUX_8525_inst
    IMB41_8526 <= IMA83_7750 when (BITSEL_u8_u1_8522_wire(0) /=  '0') else IMA82_7740;
    -- logger for split-operator MUX_8533_inst flow-through 
    process(IMB42_8534) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8533_inst:flowthrough inputs: " & " BITSEL_u8_u1_8530_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8530_wire) & " IMA85_7770 = "& Convert_SLV_To_Hex_String(IMA85_7770) & " IMA84_7760 = "& Convert_SLV_To_Hex_String(IMA84_7760) & " outputs:" & " IMB42_8534= "  & Convert_SLV_To_Hex_String(IMB42_8534));
      --
    end process; 
    -- flow-through select operator MUX_8533_inst
    IMB42_8534 <= IMA85_7770 when (BITSEL_u8_u1_8530_wire(0) /=  '0') else IMA84_7760;
    -- logger for split-operator MUX_8541_inst flow-through 
    process(IMB43_8542) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8541_inst:flowthrough inputs: " & " BITSEL_u8_u1_8538_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8538_wire) & " IMA87_7790 = "& Convert_SLV_To_Hex_String(IMA87_7790) & " IMA86_7780 = "& Convert_SLV_To_Hex_String(IMA86_7780) & " outputs:" & " IMB43_8542= "  & Convert_SLV_To_Hex_String(IMB43_8542));
      --
    end process; 
    -- flow-through select operator MUX_8541_inst
    IMB43_8542 <= IMA87_7790 when (BITSEL_u8_u1_8538_wire(0) /=  '0') else IMA86_7780;
    -- logger for split-operator MUX_8549_inst flow-through 
    process(IMB44_8550) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8549_inst:flowthrough inputs: " & " BITSEL_u8_u1_8546_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8546_wire) & " IMA89_7810 = "& Convert_SLV_To_Hex_String(IMA89_7810) & " IMA88_7800 = "& Convert_SLV_To_Hex_String(IMA88_7800) & " outputs:" & " IMB44_8550= "  & Convert_SLV_To_Hex_String(IMB44_8550));
      --
    end process; 
    -- flow-through select operator MUX_8549_inst
    IMB44_8550 <= IMA89_7810 when (BITSEL_u8_u1_8546_wire(0) /=  '0') else IMA88_7800;
    -- logger for split-operator MUX_8557_inst flow-through 
    process(IMB45_8558) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8557_inst:flowthrough inputs: " & " BITSEL_u8_u1_8554_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8554_wire) & " IMA91_7830 = "& Convert_SLV_To_Hex_String(IMA91_7830) & " IMA90_7820 = "& Convert_SLV_To_Hex_String(IMA90_7820) & " outputs:" & " IMB45_8558= "  & Convert_SLV_To_Hex_String(IMB45_8558));
      --
    end process; 
    -- flow-through select operator MUX_8557_inst
    IMB45_8558 <= IMA91_7830 when (BITSEL_u8_u1_8554_wire(0) /=  '0') else IMA90_7820;
    -- logger for split-operator MUX_8565_inst flow-through 
    process(IMB46_8566) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8565_inst:flowthrough inputs: " & " BITSEL_u8_u1_8562_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8562_wire) & " IMA93_7850 = "& Convert_SLV_To_Hex_String(IMA93_7850) & " IMA92_7840 = "& Convert_SLV_To_Hex_String(IMA92_7840) & " outputs:" & " IMB46_8566= "  & Convert_SLV_To_Hex_String(IMB46_8566));
      --
    end process; 
    -- flow-through select operator MUX_8565_inst
    IMB46_8566 <= IMA93_7850 when (BITSEL_u8_u1_8562_wire(0) /=  '0') else IMA92_7840;
    -- logger for split-operator MUX_8573_inst flow-through 
    process(IMB47_8574) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8573_inst:flowthrough inputs: " & " BITSEL_u8_u1_8570_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8570_wire) & " IMA95_7870 = "& Convert_SLV_To_Hex_String(IMA95_7870) & " IMA94_7860 = "& Convert_SLV_To_Hex_String(IMA94_7860) & " outputs:" & " IMB47_8574= "  & Convert_SLV_To_Hex_String(IMB47_8574));
      --
    end process; 
    -- flow-through select operator MUX_8573_inst
    IMB47_8574 <= IMA95_7870 when (BITSEL_u8_u1_8570_wire(0) /=  '0') else IMA94_7860;
    -- logger for split-operator MUX_8581_inst flow-through 
    process(IMB48_8582) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8581_inst:flowthrough inputs: " & " BITSEL_u8_u1_8578_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8578_wire) & " IMA97_7890 = "& Convert_SLV_To_Hex_String(IMA97_7890) & " IMA96_7880 = "& Convert_SLV_To_Hex_String(IMA96_7880) & " outputs:" & " IMB48_8582= "  & Convert_SLV_To_Hex_String(IMB48_8582));
      --
    end process; 
    -- flow-through select operator MUX_8581_inst
    IMB48_8582 <= IMA97_7890 when (BITSEL_u8_u1_8578_wire(0) /=  '0') else IMA96_7880;
    -- logger for split-operator MUX_8589_inst flow-through 
    process(IMB49_8590) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8589_inst:flowthrough inputs: " & " BITSEL_u8_u1_8586_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8586_wire) & " IMA99_7910 = "& Convert_SLV_To_Hex_String(IMA99_7910) & " IMA98_7900 = "& Convert_SLV_To_Hex_String(IMA98_7900) & " outputs:" & " IMB49_8590= "  & Convert_SLV_To_Hex_String(IMB49_8590));
      --
    end process; 
    -- flow-through select operator MUX_8589_inst
    IMB49_8590 <= IMA99_7910 when (BITSEL_u8_u1_8586_wire(0) /=  '0') else IMA98_7900;
    -- logger for split-operator MUX_8597_inst flow-through 
    process(IMB50_8598) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8597_inst:flowthrough inputs: " & " BITSEL_u8_u1_8594_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8594_wire) & " IMA101_7930 = "& Convert_SLV_To_Hex_String(IMA101_7930) & " IMA100_7920 = "& Convert_SLV_To_Hex_String(IMA100_7920) & " outputs:" & " IMB50_8598= "  & Convert_SLV_To_Hex_String(IMB50_8598));
      --
    end process; 
    -- flow-through select operator MUX_8597_inst
    IMB50_8598 <= IMA101_7930 when (BITSEL_u8_u1_8594_wire(0) /=  '0') else IMA100_7920;
    -- logger for split-operator MUX_8605_inst flow-through 
    process(IMB51_8606) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8605_inst:flowthrough inputs: " & " BITSEL_u8_u1_8602_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8602_wire) & " IMA103_7950 = "& Convert_SLV_To_Hex_String(IMA103_7950) & " IMA102_7940 = "& Convert_SLV_To_Hex_String(IMA102_7940) & " outputs:" & " IMB51_8606= "  & Convert_SLV_To_Hex_String(IMB51_8606));
      --
    end process; 
    -- flow-through select operator MUX_8605_inst
    IMB51_8606 <= IMA103_7950 when (BITSEL_u8_u1_8602_wire(0) /=  '0') else IMA102_7940;
    -- logger for split-operator MUX_8613_inst flow-through 
    process(IMB52_8614) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8613_inst:flowthrough inputs: " & " BITSEL_u8_u1_8610_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8610_wire) & " IMA105_7970 = "& Convert_SLV_To_Hex_String(IMA105_7970) & " IMA104_7960 = "& Convert_SLV_To_Hex_String(IMA104_7960) & " outputs:" & " IMB52_8614= "  & Convert_SLV_To_Hex_String(IMB52_8614));
      --
    end process; 
    -- flow-through select operator MUX_8613_inst
    IMB52_8614 <= IMA105_7970 when (BITSEL_u8_u1_8610_wire(0) /=  '0') else IMA104_7960;
    -- logger for split-operator MUX_8621_inst flow-through 
    process(IMB53_8622) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8621_inst:flowthrough inputs: " & " BITSEL_u8_u1_8618_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8618_wire) & " IMA107_7990 = "& Convert_SLV_To_Hex_String(IMA107_7990) & " IMA106_7980 = "& Convert_SLV_To_Hex_String(IMA106_7980) & " outputs:" & " IMB53_8622= "  & Convert_SLV_To_Hex_String(IMB53_8622));
      --
    end process; 
    -- flow-through select operator MUX_8621_inst
    IMB53_8622 <= IMA107_7990 when (BITSEL_u8_u1_8618_wire(0) /=  '0') else IMA106_7980;
    -- logger for split-operator MUX_8629_inst flow-through 
    process(IMB54_8630) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8629_inst:flowthrough inputs: " & " BITSEL_u8_u1_8626_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8626_wire) & " IMA109_8010 = "& Convert_SLV_To_Hex_String(IMA109_8010) & " IMA108_8000 = "& Convert_SLV_To_Hex_String(IMA108_8000) & " outputs:" & " IMB54_8630= "  & Convert_SLV_To_Hex_String(IMB54_8630));
      --
    end process; 
    -- flow-through select operator MUX_8629_inst
    IMB54_8630 <= IMA109_8010 when (BITSEL_u8_u1_8626_wire(0) /=  '0') else IMA108_8000;
    -- logger for split-operator MUX_8637_inst flow-through 
    process(IMB55_8638) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8637_inst:flowthrough inputs: " & " BITSEL_u8_u1_8634_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8634_wire) & " IMA111_8030 = "& Convert_SLV_To_Hex_String(IMA111_8030) & " IMA110_8020 = "& Convert_SLV_To_Hex_String(IMA110_8020) & " outputs:" & " IMB55_8638= "  & Convert_SLV_To_Hex_String(IMB55_8638));
      --
    end process; 
    -- flow-through select operator MUX_8637_inst
    IMB55_8638 <= IMA111_8030 when (BITSEL_u8_u1_8634_wire(0) /=  '0') else IMA110_8020;
    -- logger for split-operator MUX_8645_inst flow-through 
    process(IMB56_8646) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8645_inst:flowthrough inputs: " & " BITSEL_u8_u1_8642_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8642_wire) & " IMA113_8050 = "& Convert_SLV_To_Hex_String(IMA113_8050) & " IMA112_8040 = "& Convert_SLV_To_Hex_String(IMA112_8040) & " outputs:" & " IMB56_8646= "  & Convert_SLV_To_Hex_String(IMB56_8646));
      --
    end process; 
    -- flow-through select operator MUX_8645_inst
    IMB56_8646 <= IMA113_8050 when (BITSEL_u8_u1_8642_wire(0) /=  '0') else IMA112_8040;
    -- logger for split-operator MUX_8653_inst flow-through 
    process(IMB57_8654) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8653_inst:flowthrough inputs: " & " BITSEL_u8_u1_8650_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8650_wire) & " IMA115_8070 = "& Convert_SLV_To_Hex_String(IMA115_8070) & " IMA114_8060 = "& Convert_SLV_To_Hex_String(IMA114_8060) & " outputs:" & " IMB57_8654= "  & Convert_SLV_To_Hex_String(IMB57_8654));
      --
    end process; 
    -- flow-through select operator MUX_8653_inst
    IMB57_8654 <= IMA115_8070 when (BITSEL_u8_u1_8650_wire(0) /=  '0') else IMA114_8060;
    -- logger for split-operator MUX_8661_inst flow-through 
    process(IMB58_8662) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8661_inst:flowthrough inputs: " & " BITSEL_u8_u1_8658_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8658_wire) & " IMA117_8090 = "& Convert_SLV_To_Hex_String(IMA117_8090) & " IMA116_8080 = "& Convert_SLV_To_Hex_String(IMA116_8080) & " outputs:" & " IMB58_8662= "  & Convert_SLV_To_Hex_String(IMB58_8662));
      --
    end process; 
    -- flow-through select operator MUX_8661_inst
    IMB58_8662 <= IMA117_8090 when (BITSEL_u8_u1_8658_wire(0) /=  '0') else IMA116_8080;
    -- logger for split-operator MUX_8669_inst flow-through 
    process(IMB59_8670) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8669_inst:flowthrough inputs: " & " BITSEL_u8_u1_8666_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8666_wire) & " IMA119_8110 = "& Convert_SLV_To_Hex_String(IMA119_8110) & " IMA118_8100 = "& Convert_SLV_To_Hex_String(IMA118_8100) & " outputs:" & " IMB59_8670= "  & Convert_SLV_To_Hex_String(IMB59_8670));
      --
    end process; 
    -- flow-through select operator MUX_8669_inst
    IMB59_8670 <= IMA119_8110 when (BITSEL_u8_u1_8666_wire(0) /=  '0') else IMA118_8100;
    -- logger for split-operator MUX_8677_inst flow-through 
    process(IMB60_8678) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8677_inst:flowthrough inputs: " & " BITSEL_u8_u1_8674_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8674_wire) & " IMA121_8130 = "& Convert_SLV_To_Hex_String(IMA121_8130) & " IMA120_8120 = "& Convert_SLV_To_Hex_String(IMA120_8120) & " outputs:" & " IMB60_8678= "  & Convert_SLV_To_Hex_String(IMB60_8678));
      --
    end process; 
    -- flow-through select operator MUX_8677_inst
    IMB60_8678 <= IMA121_8130 when (BITSEL_u8_u1_8674_wire(0) /=  '0') else IMA120_8120;
    -- logger for split-operator MUX_8685_inst flow-through 
    process(IMB61_8686) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8685_inst:flowthrough inputs: " & " BITSEL_u8_u1_8682_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8682_wire) & " IMA123_8150 = "& Convert_SLV_To_Hex_String(IMA123_8150) & " IMA122_8140 = "& Convert_SLV_To_Hex_String(IMA122_8140) & " outputs:" & " IMB61_8686= "  & Convert_SLV_To_Hex_String(IMB61_8686));
      --
    end process; 
    -- flow-through select operator MUX_8685_inst
    IMB61_8686 <= IMA123_8150 when (BITSEL_u8_u1_8682_wire(0) /=  '0') else IMA122_8140;
    -- logger for split-operator MUX_8693_inst flow-through 
    process(IMB62_8694) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8693_inst:flowthrough inputs: " & " BITSEL_u8_u1_8690_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8690_wire) & " IMA125_8170 = "& Convert_SLV_To_Hex_String(IMA125_8170) & " IMA124_8160 = "& Convert_SLV_To_Hex_String(IMA124_8160) & " outputs:" & " IMB62_8694= "  & Convert_SLV_To_Hex_String(IMB62_8694));
      --
    end process; 
    -- flow-through select operator MUX_8693_inst
    IMB62_8694 <= IMA125_8170 when (BITSEL_u8_u1_8690_wire(0) /=  '0') else IMA124_8160;
    -- logger for split-operator MUX_8701_inst flow-through 
    process(IMB63_8702) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8701_inst:flowthrough inputs: " & " BITSEL_u8_u1_8698_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8698_wire) & " IMA127_8190 = "& Convert_SLV_To_Hex_String(IMA127_8190) & " IMA126_8180 = "& Convert_SLV_To_Hex_String(IMA126_8180) & " outputs:" & " IMB63_8702= "  & Convert_SLV_To_Hex_String(IMB63_8702));
      --
    end process; 
    -- flow-through select operator MUX_8701_inst
    IMB63_8702 <= IMA127_8190 when (BITSEL_u8_u1_8698_wire(0) /=  '0') else IMA126_8180;
    -- logger for split-operator MUX_8709_inst flow-through 
    process(IMC0_8710) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8709_inst:flowthrough inputs: " & " BITSEL_u8_u1_8706_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8706_wire) & " IMB1_8206 = "& Convert_SLV_To_Hex_String(IMB1_8206) & " IMB0_8198 = "& Convert_SLV_To_Hex_String(IMB0_8198) & " outputs:" & " IMC0_8710= "  & Convert_SLV_To_Hex_String(IMC0_8710));
      --
    end process; 
    -- flow-through select operator MUX_8709_inst
    IMC0_8710 <= IMB1_8206 when (BITSEL_u8_u1_8706_wire(0) /=  '0') else IMB0_8198;
    -- logger for split-operator MUX_8717_inst flow-through 
    process(IMC1_8718) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8717_inst:flowthrough inputs: " & " BITSEL_u8_u1_8714_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8714_wire) & " IMB3_8222 = "& Convert_SLV_To_Hex_String(IMB3_8222) & " IMB2_8214 = "& Convert_SLV_To_Hex_String(IMB2_8214) & " outputs:" & " IMC1_8718= "  & Convert_SLV_To_Hex_String(IMC1_8718));
      --
    end process; 
    -- flow-through select operator MUX_8717_inst
    IMC1_8718 <= IMB3_8222 when (BITSEL_u8_u1_8714_wire(0) /=  '0') else IMB2_8214;
    -- logger for split-operator MUX_8725_inst flow-through 
    process(IMC2_8726) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8725_inst:flowthrough inputs: " & " BITSEL_u8_u1_8722_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8722_wire) & " IMB5_8238 = "& Convert_SLV_To_Hex_String(IMB5_8238) & " IMB4_8230 = "& Convert_SLV_To_Hex_String(IMB4_8230) & " outputs:" & " IMC2_8726= "  & Convert_SLV_To_Hex_String(IMC2_8726));
      --
    end process; 
    -- flow-through select operator MUX_8725_inst
    IMC2_8726 <= IMB5_8238 when (BITSEL_u8_u1_8722_wire(0) /=  '0') else IMB4_8230;
    -- logger for split-operator MUX_8733_inst flow-through 
    process(IMC3_8734) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8733_inst:flowthrough inputs: " & " BITSEL_u8_u1_8730_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8730_wire) & " IMB7_8254 = "& Convert_SLV_To_Hex_String(IMB7_8254) & " IMB6_8246 = "& Convert_SLV_To_Hex_String(IMB6_8246) & " outputs:" & " IMC3_8734= "  & Convert_SLV_To_Hex_String(IMC3_8734));
      --
    end process; 
    -- flow-through select operator MUX_8733_inst
    IMC3_8734 <= IMB7_8254 when (BITSEL_u8_u1_8730_wire(0) /=  '0') else IMB6_8246;
    -- logger for split-operator MUX_8741_inst flow-through 
    process(IMC4_8742) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8741_inst:flowthrough inputs: " & " BITSEL_u8_u1_8738_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8738_wire) & " IMB9_8270 = "& Convert_SLV_To_Hex_String(IMB9_8270) & " IMB8_8262 = "& Convert_SLV_To_Hex_String(IMB8_8262) & " outputs:" & " IMC4_8742= "  & Convert_SLV_To_Hex_String(IMC4_8742));
      --
    end process; 
    -- flow-through select operator MUX_8741_inst
    IMC4_8742 <= IMB9_8270 when (BITSEL_u8_u1_8738_wire(0) /=  '0') else IMB8_8262;
    -- logger for split-operator MUX_8749_inst flow-through 
    process(IMC5_8750) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8749_inst:flowthrough inputs: " & " BITSEL_u8_u1_8746_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8746_wire) & " IMB11_8286 = "& Convert_SLV_To_Hex_String(IMB11_8286) & " IMB10_8278 = "& Convert_SLV_To_Hex_String(IMB10_8278) & " outputs:" & " IMC5_8750= "  & Convert_SLV_To_Hex_String(IMC5_8750));
      --
    end process; 
    -- flow-through select operator MUX_8749_inst
    IMC5_8750 <= IMB11_8286 when (BITSEL_u8_u1_8746_wire(0) /=  '0') else IMB10_8278;
    -- logger for split-operator MUX_8757_inst flow-through 
    process(IMC6_8758) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8757_inst:flowthrough inputs: " & " BITSEL_u8_u1_8754_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8754_wire) & " IMB13_8302 = "& Convert_SLV_To_Hex_String(IMB13_8302) & " IMB12_8294 = "& Convert_SLV_To_Hex_String(IMB12_8294) & " outputs:" & " IMC6_8758= "  & Convert_SLV_To_Hex_String(IMC6_8758));
      --
    end process; 
    -- flow-through select operator MUX_8757_inst
    IMC6_8758 <= IMB13_8302 when (BITSEL_u8_u1_8754_wire(0) /=  '0') else IMB12_8294;
    -- logger for split-operator MUX_8765_inst flow-through 
    process(IMC7_8766) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8765_inst:flowthrough inputs: " & " BITSEL_u8_u1_8762_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8762_wire) & " IMB15_8318 = "& Convert_SLV_To_Hex_String(IMB15_8318) & " IMB14_8310 = "& Convert_SLV_To_Hex_String(IMB14_8310) & " outputs:" & " IMC7_8766= "  & Convert_SLV_To_Hex_String(IMC7_8766));
      --
    end process; 
    -- flow-through select operator MUX_8765_inst
    IMC7_8766 <= IMB15_8318 when (BITSEL_u8_u1_8762_wire(0) /=  '0') else IMB14_8310;
    -- logger for split-operator MUX_8773_inst flow-through 
    process(IMC8_8774) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8773_inst:flowthrough inputs: " & " BITSEL_u8_u1_8770_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8770_wire) & " IMB17_8334 = "& Convert_SLV_To_Hex_String(IMB17_8334) & " IMB16_8326 = "& Convert_SLV_To_Hex_String(IMB16_8326) & " outputs:" & " IMC8_8774= "  & Convert_SLV_To_Hex_String(IMC8_8774));
      --
    end process; 
    -- flow-through select operator MUX_8773_inst
    IMC8_8774 <= IMB17_8334 when (BITSEL_u8_u1_8770_wire(0) /=  '0') else IMB16_8326;
    -- logger for split-operator MUX_8781_inst flow-through 
    process(IMC9_8782) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8781_inst:flowthrough inputs: " & " BITSEL_u8_u1_8778_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8778_wire) & " IMB19_8350 = "& Convert_SLV_To_Hex_String(IMB19_8350) & " IMB18_8342 = "& Convert_SLV_To_Hex_String(IMB18_8342) & " outputs:" & " IMC9_8782= "  & Convert_SLV_To_Hex_String(IMC9_8782));
      --
    end process; 
    -- flow-through select operator MUX_8781_inst
    IMC9_8782 <= IMB19_8350 when (BITSEL_u8_u1_8778_wire(0) /=  '0') else IMB18_8342;
    -- logger for split-operator MUX_8789_inst flow-through 
    process(IMC10_8790) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8789_inst:flowthrough inputs: " & " BITSEL_u8_u1_8786_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8786_wire) & " IMB21_8366 = "& Convert_SLV_To_Hex_String(IMB21_8366) & " IMB20_8358 = "& Convert_SLV_To_Hex_String(IMB20_8358) & " outputs:" & " IMC10_8790= "  & Convert_SLV_To_Hex_String(IMC10_8790));
      --
    end process; 
    -- flow-through select operator MUX_8789_inst
    IMC10_8790 <= IMB21_8366 when (BITSEL_u8_u1_8786_wire(0) /=  '0') else IMB20_8358;
    -- logger for split-operator MUX_8797_inst flow-through 
    process(IMC11_8798) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8797_inst:flowthrough inputs: " & " BITSEL_u8_u1_8794_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8794_wire) & " IMB23_8382 = "& Convert_SLV_To_Hex_String(IMB23_8382) & " IMB22_8374 = "& Convert_SLV_To_Hex_String(IMB22_8374) & " outputs:" & " IMC11_8798= "  & Convert_SLV_To_Hex_String(IMC11_8798));
      --
    end process; 
    -- flow-through select operator MUX_8797_inst
    IMC11_8798 <= IMB23_8382 when (BITSEL_u8_u1_8794_wire(0) /=  '0') else IMB22_8374;
    -- logger for split-operator MUX_8805_inst flow-through 
    process(IMC12_8806) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8805_inst:flowthrough inputs: " & " BITSEL_u8_u1_8802_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8802_wire) & " IMB25_8398 = "& Convert_SLV_To_Hex_String(IMB25_8398) & " IMB24_8390 = "& Convert_SLV_To_Hex_String(IMB24_8390) & " outputs:" & " IMC12_8806= "  & Convert_SLV_To_Hex_String(IMC12_8806));
      --
    end process; 
    -- flow-through select operator MUX_8805_inst
    IMC12_8806 <= IMB25_8398 when (BITSEL_u8_u1_8802_wire(0) /=  '0') else IMB24_8390;
    -- logger for split-operator MUX_8813_inst flow-through 
    process(IMC13_8814) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8813_inst:flowthrough inputs: " & " BITSEL_u8_u1_8810_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8810_wire) & " IMB27_8414 = "& Convert_SLV_To_Hex_String(IMB27_8414) & " IMB26_8406 = "& Convert_SLV_To_Hex_String(IMB26_8406) & " outputs:" & " IMC13_8814= "  & Convert_SLV_To_Hex_String(IMC13_8814));
      --
    end process; 
    -- flow-through select operator MUX_8813_inst
    IMC13_8814 <= IMB27_8414 when (BITSEL_u8_u1_8810_wire(0) /=  '0') else IMB26_8406;
    -- logger for split-operator MUX_8821_inst flow-through 
    process(IMC14_8822) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8821_inst:flowthrough inputs: " & " BITSEL_u8_u1_8818_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8818_wire) & " IMB29_8430 = "& Convert_SLV_To_Hex_String(IMB29_8430) & " IMB28_8422 = "& Convert_SLV_To_Hex_String(IMB28_8422) & " outputs:" & " IMC14_8822= "  & Convert_SLV_To_Hex_String(IMC14_8822));
      --
    end process; 
    -- flow-through select operator MUX_8821_inst
    IMC14_8822 <= IMB29_8430 when (BITSEL_u8_u1_8818_wire(0) /=  '0') else IMB28_8422;
    -- logger for split-operator MUX_8829_inst flow-through 
    process(IMC15_8830) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8829_inst:flowthrough inputs: " & " BITSEL_u8_u1_8826_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8826_wire) & " IMB31_8446 = "& Convert_SLV_To_Hex_String(IMB31_8446) & " IMB30_8438 = "& Convert_SLV_To_Hex_String(IMB30_8438) & " outputs:" & " IMC15_8830= "  & Convert_SLV_To_Hex_String(IMC15_8830));
      --
    end process; 
    -- flow-through select operator MUX_8829_inst
    IMC15_8830 <= IMB31_8446 when (BITSEL_u8_u1_8826_wire(0) /=  '0') else IMB30_8438;
    -- logger for split-operator MUX_8837_inst flow-through 
    process(IMC16_8838) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8837_inst:flowthrough inputs: " & " BITSEL_u8_u1_8834_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8834_wire) & " IMB33_8462 = "& Convert_SLV_To_Hex_String(IMB33_8462) & " IMB32_8454 = "& Convert_SLV_To_Hex_String(IMB32_8454) & " outputs:" & " IMC16_8838= "  & Convert_SLV_To_Hex_String(IMC16_8838));
      --
    end process; 
    -- flow-through select operator MUX_8837_inst
    IMC16_8838 <= IMB33_8462 when (BITSEL_u8_u1_8834_wire(0) /=  '0') else IMB32_8454;
    -- logger for split-operator MUX_8845_inst flow-through 
    process(IMC17_8846) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8845_inst:flowthrough inputs: " & " BITSEL_u8_u1_8842_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8842_wire) & " IMB35_8478 = "& Convert_SLV_To_Hex_String(IMB35_8478) & " IMB34_8470 = "& Convert_SLV_To_Hex_String(IMB34_8470) & " outputs:" & " IMC17_8846= "  & Convert_SLV_To_Hex_String(IMC17_8846));
      --
    end process; 
    -- flow-through select operator MUX_8845_inst
    IMC17_8846 <= IMB35_8478 when (BITSEL_u8_u1_8842_wire(0) /=  '0') else IMB34_8470;
    -- logger for split-operator MUX_8853_inst flow-through 
    process(IMC18_8854) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8853_inst:flowthrough inputs: " & " BITSEL_u8_u1_8850_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8850_wire) & " IMB37_8494 = "& Convert_SLV_To_Hex_String(IMB37_8494) & " IMB36_8486 = "& Convert_SLV_To_Hex_String(IMB36_8486) & " outputs:" & " IMC18_8854= "  & Convert_SLV_To_Hex_String(IMC18_8854));
      --
    end process; 
    -- flow-through select operator MUX_8853_inst
    IMC18_8854 <= IMB37_8494 when (BITSEL_u8_u1_8850_wire(0) /=  '0') else IMB36_8486;
    -- logger for split-operator MUX_8861_inst flow-through 
    process(IMC19_8862) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8861_inst:flowthrough inputs: " & " BITSEL_u8_u1_8858_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8858_wire) & " IMB39_8510 = "& Convert_SLV_To_Hex_String(IMB39_8510) & " IMB38_8502 = "& Convert_SLV_To_Hex_String(IMB38_8502) & " outputs:" & " IMC19_8862= "  & Convert_SLV_To_Hex_String(IMC19_8862));
      --
    end process; 
    -- flow-through select operator MUX_8861_inst
    IMC19_8862 <= IMB39_8510 when (BITSEL_u8_u1_8858_wire(0) /=  '0') else IMB38_8502;
    -- logger for split-operator MUX_8869_inst flow-through 
    process(IMC20_8870) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8869_inst:flowthrough inputs: " & " BITSEL_u8_u1_8866_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8866_wire) & " IMB41_8526 = "& Convert_SLV_To_Hex_String(IMB41_8526) & " IMB40_8518 = "& Convert_SLV_To_Hex_String(IMB40_8518) & " outputs:" & " IMC20_8870= "  & Convert_SLV_To_Hex_String(IMC20_8870));
      --
    end process; 
    -- flow-through select operator MUX_8869_inst
    IMC20_8870 <= IMB41_8526 when (BITSEL_u8_u1_8866_wire(0) /=  '0') else IMB40_8518;
    -- logger for split-operator MUX_8877_inst flow-through 
    process(IMC21_8878) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8877_inst:flowthrough inputs: " & " BITSEL_u8_u1_8874_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8874_wire) & " IMB43_8542 = "& Convert_SLV_To_Hex_String(IMB43_8542) & " IMB42_8534 = "& Convert_SLV_To_Hex_String(IMB42_8534) & " outputs:" & " IMC21_8878= "  & Convert_SLV_To_Hex_String(IMC21_8878));
      --
    end process; 
    -- flow-through select operator MUX_8877_inst
    IMC21_8878 <= IMB43_8542 when (BITSEL_u8_u1_8874_wire(0) /=  '0') else IMB42_8534;
    -- logger for split-operator MUX_8885_inst flow-through 
    process(IMC22_8886) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8885_inst:flowthrough inputs: " & " BITSEL_u8_u1_8882_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8882_wire) & " IMB45_8558 = "& Convert_SLV_To_Hex_String(IMB45_8558) & " IMB44_8550 = "& Convert_SLV_To_Hex_String(IMB44_8550) & " outputs:" & " IMC22_8886= "  & Convert_SLV_To_Hex_String(IMC22_8886));
      --
    end process; 
    -- flow-through select operator MUX_8885_inst
    IMC22_8886 <= IMB45_8558 when (BITSEL_u8_u1_8882_wire(0) /=  '0') else IMB44_8550;
    -- logger for split-operator MUX_8893_inst flow-through 
    process(IMC23_8894) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8893_inst:flowthrough inputs: " & " BITSEL_u8_u1_8890_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8890_wire) & " IMB47_8574 = "& Convert_SLV_To_Hex_String(IMB47_8574) & " IMB46_8566 = "& Convert_SLV_To_Hex_String(IMB46_8566) & " outputs:" & " IMC23_8894= "  & Convert_SLV_To_Hex_String(IMC23_8894));
      --
    end process; 
    -- flow-through select operator MUX_8893_inst
    IMC23_8894 <= IMB47_8574 when (BITSEL_u8_u1_8890_wire(0) /=  '0') else IMB46_8566;
    -- logger for split-operator MUX_8901_inst flow-through 
    process(IMC24_8902) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8901_inst:flowthrough inputs: " & " BITSEL_u8_u1_8898_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8898_wire) & " IMB49_8590 = "& Convert_SLV_To_Hex_String(IMB49_8590) & " IMB48_8582 = "& Convert_SLV_To_Hex_String(IMB48_8582) & " outputs:" & " IMC24_8902= "  & Convert_SLV_To_Hex_String(IMC24_8902));
      --
    end process; 
    -- flow-through select operator MUX_8901_inst
    IMC24_8902 <= IMB49_8590 when (BITSEL_u8_u1_8898_wire(0) /=  '0') else IMB48_8582;
    -- logger for split-operator MUX_8909_inst flow-through 
    process(IMC25_8910) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8909_inst:flowthrough inputs: " & " BITSEL_u8_u1_8906_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8906_wire) & " IMB51_8606 = "& Convert_SLV_To_Hex_String(IMB51_8606) & " IMB50_8598 = "& Convert_SLV_To_Hex_String(IMB50_8598) & " outputs:" & " IMC25_8910= "  & Convert_SLV_To_Hex_String(IMC25_8910));
      --
    end process; 
    -- flow-through select operator MUX_8909_inst
    IMC25_8910 <= IMB51_8606 when (BITSEL_u8_u1_8906_wire(0) /=  '0') else IMB50_8598;
    -- logger for split-operator MUX_8917_inst flow-through 
    process(IMC26_8918) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8917_inst:flowthrough inputs: " & " BITSEL_u8_u1_8914_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8914_wire) & " IMB53_8622 = "& Convert_SLV_To_Hex_String(IMB53_8622) & " IMB52_8614 = "& Convert_SLV_To_Hex_String(IMB52_8614) & " outputs:" & " IMC26_8918= "  & Convert_SLV_To_Hex_String(IMC26_8918));
      --
    end process; 
    -- flow-through select operator MUX_8917_inst
    IMC26_8918 <= IMB53_8622 when (BITSEL_u8_u1_8914_wire(0) /=  '0') else IMB52_8614;
    -- logger for split-operator MUX_8925_inst flow-through 
    process(IMC27_8926) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8925_inst:flowthrough inputs: " & " BITSEL_u8_u1_8922_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8922_wire) & " IMB55_8638 = "& Convert_SLV_To_Hex_String(IMB55_8638) & " IMB54_8630 = "& Convert_SLV_To_Hex_String(IMB54_8630) & " outputs:" & " IMC27_8926= "  & Convert_SLV_To_Hex_String(IMC27_8926));
      --
    end process; 
    -- flow-through select operator MUX_8925_inst
    IMC27_8926 <= IMB55_8638 when (BITSEL_u8_u1_8922_wire(0) /=  '0') else IMB54_8630;
    -- logger for split-operator MUX_8933_inst flow-through 
    process(IMC28_8934) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8933_inst:flowthrough inputs: " & " BITSEL_u8_u1_8930_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8930_wire) & " IMB57_8654 = "& Convert_SLV_To_Hex_String(IMB57_8654) & " IMB56_8646 = "& Convert_SLV_To_Hex_String(IMB56_8646) & " outputs:" & " IMC28_8934= "  & Convert_SLV_To_Hex_String(IMC28_8934));
      --
    end process; 
    -- flow-through select operator MUX_8933_inst
    IMC28_8934 <= IMB57_8654 when (BITSEL_u8_u1_8930_wire(0) /=  '0') else IMB56_8646;
    -- logger for split-operator MUX_8941_inst flow-through 
    process(IMC29_8942) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8941_inst:flowthrough inputs: " & " BITSEL_u8_u1_8938_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8938_wire) & " IMB59_8670 = "& Convert_SLV_To_Hex_String(IMB59_8670) & " IMB58_8662 = "& Convert_SLV_To_Hex_String(IMB58_8662) & " outputs:" & " IMC29_8942= "  & Convert_SLV_To_Hex_String(IMC29_8942));
      --
    end process; 
    -- flow-through select operator MUX_8941_inst
    IMC29_8942 <= IMB59_8670 when (BITSEL_u8_u1_8938_wire(0) /=  '0') else IMB58_8662;
    -- logger for split-operator MUX_8949_inst flow-through 
    process(IMC30_8950) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8949_inst:flowthrough inputs: " & " BITSEL_u8_u1_8946_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8946_wire) & " IMB61_8686 = "& Convert_SLV_To_Hex_String(IMB61_8686) & " IMB60_8678 = "& Convert_SLV_To_Hex_String(IMB60_8678) & " outputs:" & " IMC30_8950= "  & Convert_SLV_To_Hex_String(IMC30_8950));
      --
    end process; 
    -- flow-through select operator MUX_8949_inst
    IMC30_8950 <= IMB61_8686 when (BITSEL_u8_u1_8946_wire(0) /=  '0') else IMB60_8678;
    -- logger for split-operator MUX_8957_inst flow-through 
    process(IMC31_8958) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8957_inst:flowthrough inputs: " & " BITSEL_u8_u1_8954_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8954_wire) & " IMB63_8702 = "& Convert_SLV_To_Hex_String(IMB63_8702) & " IMB62_8694 = "& Convert_SLV_To_Hex_String(IMB62_8694) & " outputs:" & " IMC31_8958= "  & Convert_SLV_To_Hex_String(IMC31_8958));
      --
    end process; 
    -- flow-through select operator MUX_8957_inst
    IMC31_8958 <= IMB63_8702 when (BITSEL_u8_u1_8954_wire(0) /=  '0') else IMB62_8694;
    -- logger for split-operator MUX_8965_inst flow-through 
    process(IMD0_8966) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8965_inst:flowthrough inputs: " & " BITSEL_u8_u1_8962_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8962_wire) & " IMC1_8718 = "& Convert_SLV_To_Hex_String(IMC1_8718) & " IMC0_8710 = "& Convert_SLV_To_Hex_String(IMC0_8710) & " outputs:" & " IMD0_8966= "  & Convert_SLV_To_Hex_String(IMD0_8966));
      --
    end process; 
    -- flow-through select operator MUX_8965_inst
    IMD0_8966 <= IMC1_8718 when (BITSEL_u8_u1_8962_wire(0) /=  '0') else IMC0_8710;
    -- logger for split-operator MUX_8973_inst flow-through 
    process(IMD1_8974) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8973_inst:flowthrough inputs: " & " BITSEL_u8_u1_8970_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8970_wire) & " IMC3_8734 = "& Convert_SLV_To_Hex_String(IMC3_8734) & " IMC2_8726 = "& Convert_SLV_To_Hex_String(IMC2_8726) & " outputs:" & " IMD1_8974= "  & Convert_SLV_To_Hex_String(IMD1_8974));
      --
    end process; 
    -- flow-through select operator MUX_8973_inst
    IMD1_8974 <= IMC3_8734 when (BITSEL_u8_u1_8970_wire(0) /=  '0') else IMC2_8726;
    -- logger for split-operator MUX_8981_inst flow-through 
    process(IMD2_8982) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8981_inst:flowthrough inputs: " & " BITSEL_u8_u1_8978_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8978_wire) & " IMC5_8750 = "& Convert_SLV_To_Hex_String(IMC5_8750) & " IMC4_8742 = "& Convert_SLV_To_Hex_String(IMC4_8742) & " outputs:" & " IMD2_8982= "  & Convert_SLV_To_Hex_String(IMD2_8982));
      --
    end process; 
    -- flow-through select operator MUX_8981_inst
    IMD2_8982 <= IMC5_8750 when (BITSEL_u8_u1_8978_wire(0) /=  '0') else IMC4_8742;
    -- logger for split-operator MUX_8989_inst flow-through 
    process(IMD3_8990) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8989_inst:flowthrough inputs: " & " BITSEL_u8_u1_8986_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8986_wire) & " IMC7_8766 = "& Convert_SLV_To_Hex_String(IMC7_8766) & " IMC6_8758 = "& Convert_SLV_To_Hex_String(IMC6_8758) & " outputs:" & " IMD3_8990= "  & Convert_SLV_To_Hex_String(IMD3_8990));
      --
    end process; 
    -- flow-through select operator MUX_8989_inst
    IMD3_8990 <= IMC7_8766 when (BITSEL_u8_u1_8986_wire(0) /=  '0') else IMC6_8758;
    -- logger for split-operator MUX_8997_inst flow-through 
    process(IMD4_8998) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_8997_inst:flowthrough inputs: " & " BITSEL_u8_u1_8994_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_8994_wire) & " IMC9_8782 = "& Convert_SLV_To_Hex_String(IMC9_8782) & " IMC8_8774 = "& Convert_SLV_To_Hex_String(IMC8_8774) & " outputs:" & " IMD4_8998= "  & Convert_SLV_To_Hex_String(IMD4_8998));
      --
    end process; 
    -- flow-through select operator MUX_8997_inst
    IMD4_8998 <= IMC9_8782 when (BITSEL_u8_u1_8994_wire(0) /=  '0') else IMC8_8774;
    -- logger for split-operator MUX_9005_inst flow-through 
    process(IMD5_9006) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_9005_inst:flowthrough inputs: " & " BITSEL_u8_u1_9002_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_9002_wire) & " IMC11_8798 = "& Convert_SLV_To_Hex_String(IMC11_8798) & " IMC10_8790 = "& Convert_SLV_To_Hex_String(IMC10_8790) & " outputs:" & " IMD5_9006= "  & Convert_SLV_To_Hex_String(IMD5_9006));
      --
    end process; 
    -- flow-through select operator MUX_9005_inst
    IMD5_9006 <= IMC11_8798 when (BITSEL_u8_u1_9002_wire(0) /=  '0') else IMC10_8790;
    -- logger for split-operator MUX_9013_inst flow-through 
    process(IMD6_9014) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_9013_inst:flowthrough inputs: " & " BITSEL_u8_u1_9010_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_9010_wire) & " IMC13_8814 = "& Convert_SLV_To_Hex_String(IMC13_8814) & " IMC12_8806 = "& Convert_SLV_To_Hex_String(IMC12_8806) & " outputs:" & " IMD6_9014= "  & Convert_SLV_To_Hex_String(IMD6_9014));
      --
    end process; 
    -- flow-through select operator MUX_9013_inst
    IMD6_9014 <= IMC13_8814 when (BITSEL_u8_u1_9010_wire(0) /=  '0') else IMC12_8806;
    -- logger for split-operator MUX_9021_inst flow-through 
    process(IMD7_9022) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_9021_inst:flowthrough inputs: " & " BITSEL_u8_u1_9018_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_9018_wire) & " IMC15_8830 = "& Convert_SLV_To_Hex_String(IMC15_8830) & " IMC14_8822 = "& Convert_SLV_To_Hex_String(IMC14_8822) & " outputs:" & " IMD7_9022= "  & Convert_SLV_To_Hex_String(IMD7_9022));
      --
    end process; 
    -- flow-through select operator MUX_9021_inst
    IMD7_9022 <= IMC15_8830 when (BITSEL_u8_u1_9018_wire(0) /=  '0') else IMC14_8822;
    -- logger for split-operator MUX_9029_inst flow-through 
    process(IMD8_9030) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_9029_inst:flowthrough inputs: " & " BITSEL_u8_u1_9026_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_9026_wire) & " IMC17_8846 = "& Convert_SLV_To_Hex_String(IMC17_8846) & " IMC16_8838 = "& Convert_SLV_To_Hex_String(IMC16_8838) & " outputs:" & " IMD8_9030= "  & Convert_SLV_To_Hex_String(IMD8_9030));
      --
    end process; 
    -- flow-through select operator MUX_9029_inst
    IMD8_9030 <= IMC17_8846 when (BITSEL_u8_u1_9026_wire(0) /=  '0') else IMC16_8838;
    -- logger for split-operator MUX_9037_inst flow-through 
    process(IMD9_9038) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_9037_inst:flowthrough inputs: " & " BITSEL_u8_u1_9034_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_9034_wire) & " IMC19_8862 = "& Convert_SLV_To_Hex_String(IMC19_8862) & " IMC18_8854 = "& Convert_SLV_To_Hex_String(IMC18_8854) & " outputs:" & " IMD9_9038= "  & Convert_SLV_To_Hex_String(IMD9_9038));
      --
    end process; 
    -- flow-through select operator MUX_9037_inst
    IMD9_9038 <= IMC19_8862 when (BITSEL_u8_u1_9034_wire(0) /=  '0') else IMC18_8854;
    -- logger for split-operator MUX_9045_inst flow-through 
    process(IMD10_9046) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_9045_inst:flowthrough inputs: " & " BITSEL_u8_u1_9042_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_9042_wire) & " IMC21_8878 = "& Convert_SLV_To_Hex_String(IMC21_8878) & " IMC20_8870 = "& Convert_SLV_To_Hex_String(IMC20_8870) & " outputs:" & " IMD10_9046= "  & Convert_SLV_To_Hex_String(IMD10_9046));
      --
    end process; 
    -- flow-through select operator MUX_9045_inst
    IMD10_9046 <= IMC21_8878 when (BITSEL_u8_u1_9042_wire(0) /=  '0') else IMC20_8870;
    -- logger for split-operator MUX_9053_inst flow-through 
    process(IMD11_9054) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_9053_inst:flowthrough inputs: " & " BITSEL_u8_u1_9050_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_9050_wire) & " IMC23_8894 = "& Convert_SLV_To_Hex_String(IMC23_8894) & " IMC22_8886 = "& Convert_SLV_To_Hex_String(IMC22_8886) & " outputs:" & " IMD11_9054= "  & Convert_SLV_To_Hex_String(IMD11_9054));
      --
    end process; 
    -- flow-through select operator MUX_9053_inst
    IMD11_9054 <= IMC23_8894 when (BITSEL_u8_u1_9050_wire(0) /=  '0') else IMC22_8886;
    -- logger for split-operator MUX_9061_inst flow-through 
    process(IMD12_9062) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_9061_inst:flowthrough inputs: " & " BITSEL_u8_u1_9058_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_9058_wire) & " IMC25_8910 = "& Convert_SLV_To_Hex_String(IMC25_8910) & " IMC24_8902 = "& Convert_SLV_To_Hex_String(IMC24_8902) & " outputs:" & " IMD12_9062= "  & Convert_SLV_To_Hex_String(IMD12_9062));
      --
    end process; 
    -- flow-through select operator MUX_9061_inst
    IMD12_9062 <= IMC25_8910 when (BITSEL_u8_u1_9058_wire(0) /=  '0') else IMC24_8902;
    -- logger for split-operator MUX_9069_inst flow-through 
    process(IMD13_9070) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_9069_inst:flowthrough inputs: " & " BITSEL_u8_u1_9066_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_9066_wire) & " IMC27_8926 = "& Convert_SLV_To_Hex_String(IMC27_8926) & " IMC26_8918 = "& Convert_SLV_To_Hex_String(IMC26_8918) & " outputs:" & " IMD13_9070= "  & Convert_SLV_To_Hex_String(IMD13_9070));
      --
    end process; 
    -- flow-through select operator MUX_9069_inst
    IMD13_9070 <= IMC27_8926 when (BITSEL_u8_u1_9066_wire(0) /=  '0') else IMC26_8918;
    -- logger for split-operator MUX_9077_inst flow-through 
    process(IMD14_9078) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_9077_inst:flowthrough inputs: " & " BITSEL_u8_u1_9074_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_9074_wire) & " IMC29_8942 = "& Convert_SLV_To_Hex_String(IMC29_8942) & " IMC28_8934 = "& Convert_SLV_To_Hex_String(IMC28_8934) & " outputs:" & " IMD14_9078= "  & Convert_SLV_To_Hex_String(IMD14_9078));
      --
    end process; 
    -- flow-through select operator MUX_9077_inst
    IMD14_9078 <= IMC29_8942 when (BITSEL_u8_u1_9074_wire(0) /=  '0') else IMC28_8934;
    -- logger for split-operator MUX_9085_inst flow-through 
    process(IMD15_9086) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_9085_inst:flowthrough inputs: " & " BITSEL_u8_u1_9082_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_9082_wire) & " IMC31_8958 = "& Convert_SLV_To_Hex_String(IMC31_8958) & " IMC30_8950 = "& Convert_SLV_To_Hex_String(IMC30_8950) & " outputs:" & " IMD15_9086= "  & Convert_SLV_To_Hex_String(IMD15_9086));
      --
    end process; 
    -- flow-through select operator MUX_9085_inst
    IMD15_9086 <= IMC31_8958 when (BITSEL_u8_u1_9082_wire(0) /=  '0') else IMC30_8950;
    -- logger for split-operator MUX_9093_inst flow-through 
    process(IME0_9094) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_9093_inst:flowthrough inputs: " & " BITSEL_u8_u1_9090_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_9090_wire) & " IMD1_8974 = "& Convert_SLV_To_Hex_String(IMD1_8974) & " IMD0_8966 = "& Convert_SLV_To_Hex_String(IMD0_8966) & " outputs:" & " IME0_9094= "  & Convert_SLV_To_Hex_String(IME0_9094));
      --
    end process; 
    -- flow-through select operator MUX_9093_inst
    IME0_9094 <= IMD1_8974 when (BITSEL_u8_u1_9090_wire(0) /=  '0') else IMD0_8966;
    -- logger for split-operator MUX_9101_inst flow-through 
    process(IME1_9102) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_9101_inst:flowthrough inputs: " & " BITSEL_u8_u1_9098_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_9098_wire) & " IMD3_8990 = "& Convert_SLV_To_Hex_String(IMD3_8990) & " IMD2_8982 = "& Convert_SLV_To_Hex_String(IMD2_8982) & " outputs:" & " IME1_9102= "  & Convert_SLV_To_Hex_String(IME1_9102));
      --
    end process; 
    -- flow-through select operator MUX_9101_inst
    IME1_9102 <= IMD3_8990 when (BITSEL_u8_u1_9098_wire(0) /=  '0') else IMD2_8982;
    -- logger for split-operator MUX_9109_inst flow-through 
    process(IME2_9110) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_9109_inst:flowthrough inputs: " & " BITSEL_u8_u1_9106_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_9106_wire) & " IMD5_9006 = "& Convert_SLV_To_Hex_String(IMD5_9006) & " IMD4_8998 = "& Convert_SLV_To_Hex_String(IMD4_8998) & " outputs:" & " IME2_9110= "  & Convert_SLV_To_Hex_String(IME2_9110));
      --
    end process; 
    -- flow-through select operator MUX_9109_inst
    IME2_9110 <= IMD5_9006 when (BITSEL_u8_u1_9106_wire(0) /=  '0') else IMD4_8998;
    -- logger for split-operator MUX_9117_inst flow-through 
    process(IME3_9118) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_9117_inst:flowthrough inputs: " & " BITSEL_u8_u1_9114_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_9114_wire) & " IMD7_9022 = "& Convert_SLV_To_Hex_String(IMD7_9022) & " IMD6_9014 = "& Convert_SLV_To_Hex_String(IMD6_9014) & " outputs:" & " IME3_9118= "  & Convert_SLV_To_Hex_String(IME3_9118));
      --
    end process; 
    -- flow-through select operator MUX_9117_inst
    IME3_9118 <= IMD7_9022 when (BITSEL_u8_u1_9114_wire(0) /=  '0') else IMD6_9014;
    -- logger for split-operator MUX_9125_inst flow-through 
    process(IME4_9126) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_9125_inst:flowthrough inputs: " & " BITSEL_u8_u1_9122_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_9122_wire) & " IMD9_9038 = "& Convert_SLV_To_Hex_String(IMD9_9038) & " IMD8_9030 = "& Convert_SLV_To_Hex_String(IMD8_9030) & " outputs:" & " IME4_9126= "  & Convert_SLV_To_Hex_String(IME4_9126));
      --
    end process; 
    -- flow-through select operator MUX_9125_inst
    IME4_9126 <= IMD9_9038 when (BITSEL_u8_u1_9122_wire(0) /=  '0') else IMD8_9030;
    -- logger for split-operator MUX_9133_inst flow-through 
    process(IME5_9134) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_9133_inst:flowthrough inputs: " & " BITSEL_u8_u1_9130_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_9130_wire) & " IMD11_9054 = "& Convert_SLV_To_Hex_String(IMD11_9054) & " IMD10_9046 = "& Convert_SLV_To_Hex_String(IMD10_9046) & " outputs:" & " IME5_9134= "  & Convert_SLV_To_Hex_String(IME5_9134));
      --
    end process; 
    -- flow-through select operator MUX_9133_inst
    IME5_9134 <= IMD11_9054 when (BITSEL_u8_u1_9130_wire(0) /=  '0') else IMD10_9046;
    -- logger for split-operator MUX_9141_inst flow-through 
    process(IME6_9142) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_9141_inst:flowthrough inputs: " & " BITSEL_u8_u1_9138_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_9138_wire) & " IMD13_9070 = "& Convert_SLV_To_Hex_String(IMD13_9070) & " IMD12_9062 = "& Convert_SLV_To_Hex_String(IMD12_9062) & " outputs:" & " IME6_9142= "  & Convert_SLV_To_Hex_String(IME6_9142));
      --
    end process; 
    -- flow-through select operator MUX_9141_inst
    IME6_9142 <= IMD13_9070 when (BITSEL_u8_u1_9138_wire(0) /=  '0') else IMD12_9062;
    -- logger for split-operator MUX_9149_inst flow-through 
    process(IME7_9150) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_9149_inst:flowthrough inputs: " & " BITSEL_u8_u1_9146_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_9146_wire) & " IMD15_9086 = "& Convert_SLV_To_Hex_String(IMD15_9086) & " IMD14_9078 = "& Convert_SLV_To_Hex_String(IMD14_9078) & " outputs:" & " IME7_9150= "  & Convert_SLV_To_Hex_String(IME7_9150));
      --
    end process; 
    -- flow-through select operator MUX_9149_inst
    IME7_9150 <= IMD15_9086 when (BITSEL_u8_u1_9146_wire(0) /=  '0') else IMD14_9078;
    -- logger for split-operator MUX_9157_inst flow-through 
    process(IMF0_9158) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_9157_inst:flowthrough inputs: " & " BITSEL_u8_u1_9154_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_9154_wire) & " IME1_9102 = "& Convert_SLV_To_Hex_String(IME1_9102) & " IME0_9094 = "& Convert_SLV_To_Hex_String(IME0_9094) & " outputs:" & " IMF0_9158= "  & Convert_SLV_To_Hex_String(IMF0_9158));
      --
    end process; 
    -- flow-through select operator MUX_9157_inst
    IMF0_9158 <= IME1_9102 when (BITSEL_u8_u1_9154_wire(0) /=  '0') else IME0_9094;
    -- logger for split-operator MUX_9165_inst flow-through 
    process(IMF1_9166) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_9165_inst:flowthrough inputs: " & " BITSEL_u8_u1_9162_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_9162_wire) & " IME3_9118 = "& Convert_SLV_To_Hex_String(IME3_9118) & " IME2_9110 = "& Convert_SLV_To_Hex_String(IME2_9110) & " outputs:" & " IMF1_9166= "  & Convert_SLV_To_Hex_String(IMF1_9166));
      --
    end process; 
    -- flow-through select operator MUX_9165_inst
    IMF1_9166 <= IME3_9118 when (BITSEL_u8_u1_9162_wire(0) /=  '0') else IME2_9110;
    -- logger for split-operator MUX_9173_inst flow-through 
    process(IMF2_9174) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_9173_inst:flowthrough inputs: " & " BITSEL_u8_u1_9170_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_9170_wire) & " IME5_9134 = "& Convert_SLV_To_Hex_String(IME5_9134) & " IME4_9126 = "& Convert_SLV_To_Hex_String(IME4_9126) & " outputs:" & " IMF2_9174= "  & Convert_SLV_To_Hex_String(IMF2_9174));
      --
    end process; 
    -- flow-through select operator MUX_9173_inst
    IMF2_9174 <= IME5_9134 when (BITSEL_u8_u1_9170_wire(0) /=  '0') else IME4_9126;
    -- logger for split-operator MUX_9181_inst flow-through 
    process(IMF3_9182) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_9181_inst:flowthrough inputs: " & " BITSEL_u8_u1_9178_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_9178_wire) & " IME7_9150 = "& Convert_SLV_To_Hex_String(IME7_9150) & " IME6_9142 = "& Convert_SLV_To_Hex_String(IME6_9142) & " outputs:" & " IMF3_9182= "  & Convert_SLV_To_Hex_String(IMF3_9182));
      --
    end process; 
    -- flow-through select operator MUX_9181_inst
    IMF3_9182 <= IME7_9150 when (BITSEL_u8_u1_9178_wire(0) /=  '0') else IME6_9142;
    -- logger for split-operator MUX_9189_inst flow-through 
    process(IMG0_9190) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_9189_inst:flowthrough inputs: " & " BITSEL_u8_u1_9186_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_9186_wire) & " IMF1_9166 = "& Convert_SLV_To_Hex_String(IMF1_9166) & " IMF0_9158 = "& Convert_SLV_To_Hex_String(IMF0_9158) & " outputs:" & " IMG0_9190= "  & Convert_SLV_To_Hex_String(IMG0_9190));
      --
    end process; 
    -- flow-through select operator MUX_9189_inst
    IMG0_9190 <= IMF1_9166 when (BITSEL_u8_u1_9186_wire(0) /=  '0') else IMF0_9158;
    -- logger for split-operator MUX_9197_inst flow-through 
    process(IMG1_9198) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_9197_inst:flowthrough inputs: " & " BITSEL_u8_u1_9194_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_9194_wire) & " IMF3_9182 = "& Convert_SLV_To_Hex_String(IMF3_9182) & " IMF2_9174 = "& Convert_SLV_To_Hex_String(IMF2_9174) & " outputs:" & " IMG1_9198= "  & Convert_SLV_To_Hex_String(IMG1_9198));
      --
    end process; 
    -- flow-through select operator MUX_9197_inst
    IMG1_9198 <= IMF3_9182 when (BITSEL_u8_u1_9194_wire(0) /=  '0') else IMF2_9174;
    -- logger for split-operator MUX_9205_inst flow-through 
    process(s_out_buffer) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:MUX_9205_inst:flowthrough inputs: " & " BITSEL_u8_u1_9202_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_9202_wire) & " IMG1_9198 = "& Convert_SLV_To_Hex_String(IMG1_9198) & " IMG0_9190 = "& Convert_SLV_To_Hex_String(IMG0_9190) & " outputs:" & " s_out_buffer= "  & Convert_SLV_To_Hex_String(s_out_buffer));
      --
    end process; 
    -- flow-through select operator MUX_9205_inst
    s_out_buffer <= IMG1_9198 when (BITSEL_u8_u1_9202_wire(0) /=  '0') else IMG0_9190;
    -- logger for split-operator BITSEL_u8_u1_6914_inst flow-through 
    process(BITSEL_u8_u1_6914_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_6914_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6913_wire_constant = "& Convert_SLV_To_Hex_String(konst_6913_wire_constant) & " outputs:" & " BITSEL_u8_u1_6914_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6914_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6914_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6913_wire_constant, tmp_var);
      BITSEL_u8_u1_6914_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6924_inst flow-through 
    process(BITSEL_u8_u1_6924_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_6924_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6923_wire_constant = "& Convert_SLV_To_Hex_String(konst_6923_wire_constant) & " outputs:" & " BITSEL_u8_u1_6924_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6924_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6924_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6923_wire_constant, tmp_var);
      BITSEL_u8_u1_6924_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6934_inst flow-through 
    process(BITSEL_u8_u1_6934_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_6934_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6933_wire_constant = "& Convert_SLV_To_Hex_String(konst_6933_wire_constant) & " outputs:" & " BITSEL_u8_u1_6934_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6934_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6934_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6933_wire_constant, tmp_var);
      BITSEL_u8_u1_6934_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6944_inst flow-through 
    process(BITSEL_u8_u1_6944_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_6944_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6943_wire_constant = "& Convert_SLV_To_Hex_String(konst_6943_wire_constant) & " outputs:" & " BITSEL_u8_u1_6944_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6944_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6944_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6943_wire_constant, tmp_var);
      BITSEL_u8_u1_6944_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6954_inst flow-through 
    process(BITSEL_u8_u1_6954_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_6954_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6953_wire_constant = "& Convert_SLV_To_Hex_String(konst_6953_wire_constant) & " outputs:" & " BITSEL_u8_u1_6954_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6954_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6954_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6953_wire_constant, tmp_var);
      BITSEL_u8_u1_6954_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6964_inst flow-through 
    process(BITSEL_u8_u1_6964_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_6964_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6963_wire_constant = "& Convert_SLV_To_Hex_String(konst_6963_wire_constant) & " outputs:" & " BITSEL_u8_u1_6964_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6964_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6964_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6963_wire_constant, tmp_var);
      BITSEL_u8_u1_6964_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6974_inst flow-through 
    process(BITSEL_u8_u1_6974_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_6974_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6973_wire_constant = "& Convert_SLV_To_Hex_String(konst_6973_wire_constant) & " outputs:" & " BITSEL_u8_u1_6974_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6974_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6974_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6973_wire_constant, tmp_var);
      BITSEL_u8_u1_6974_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6984_inst flow-through 
    process(BITSEL_u8_u1_6984_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_6984_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6983_wire_constant = "& Convert_SLV_To_Hex_String(konst_6983_wire_constant) & " outputs:" & " BITSEL_u8_u1_6984_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6984_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6984_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6983_wire_constant, tmp_var);
      BITSEL_u8_u1_6984_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_6994_inst flow-through 
    process(BITSEL_u8_u1_6994_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_6994_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_6993_wire_constant = "& Convert_SLV_To_Hex_String(konst_6993_wire_constant) & " outputs:" & " BITSEL_u8_u1_6994_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_6994_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_6994_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6993_wire_constant, tmp_var);
      BITSEL_u8_u1_6994_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_7004_inst flow-through 
    process(BITSEL_u8_u1_7004_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_7004_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_7003_wire_constant = "& Convert_SLV_To_Hex_String(konst_7003_wire_constant) & " outputs:" & " BITSEL_u8_u1_7004_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_7004_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_7004_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7003_wire_constant, tmp_var);
      BITSEL_u8_u1_7004_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_7014_inst flow-through 
    process(BITSEL_u8_u1_7014_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_7014_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_7013_wire_constant = "& Convert_SLV_To_Hex_String(konst_7013_wire_constant) & " outputs:" & " BITSEL_u8_u1_7014_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_7014_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_7014_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7013_wire_constant, tmp_var);
      BITSEL_u8_u1_7014_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_7024_inst flow-through 
    process(BITSEL_u8_u1_7024_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_7024_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_7023_wire_constant = "& Convert_SLV_To_Hex_String(konst_7023_wire_constant) & " outputs:" & " BITSEL_u8_u1_7024_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_7024_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_7024_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7023_wire_constant, tmp_var);
      BITSEL_u8_u1_7024_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_7034_inst flow-through 
    process(BITSEL_u8_u1_7034_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_7034_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_7033_wire_constant = "& Convert_SLV_To_Hex_String(konst_7033_wire_constant) & " outputs:" & " BITSEL_u8_u1_7034_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_7034_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_7034_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7033_wire_constant, tmp_var);
      BITSEL_u8_u1_7034_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_7044_inst flow-through 
    process(BITSEL_u8_u1_7044_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_7044_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_7043_wire_constant = "& Convert_SLV_To_Hex_String(konst_7043_wire_constant) & " outputs:" & " BITSEL_u8_u1_7044_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_7044_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_7044_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7043_wire_constant, tmp_var);
      BITSEL_u8_u1_7044_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_7054_inst flow-through 
    process(BITSEL_u8_u1_7054_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_7054_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_7053_wire_constant = "& Convert_SLV_To_Hex_String(konst_7053_wire_constant) & " outputs:" & " BITSEL_u8_u1_7054_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_7054_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_7054_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7053_wire_constant, tmp_var);
      BITSEL_u8_u1_7054_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_7064_inst flow-through 
    process(BITSEL_u8_u1_7064_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_7064_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_7063_wire_constant = "& Convert_SLV_To_Hex_String(konst_7063_wire_constant) & " outputs:" & " BITSEL_u8_u1_7064_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_7064_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_7064_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7063_wire_constant, tmp_var);
      BITSEL_u8_u1_7064_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_7074_inst flow-through 
    process(BITSEL_u8_u1_7074_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_7074_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_7073_wire_constant = "& Convert_SLV_To_Hex_String(konst_7073_wire_constant) & " outputs:" & " BITSEL_u8_u1_7074_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_7074_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_7074_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7073_wire_constant, tmp_var);
      BITSEL_u8_u1_7074_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_7084_inst flow-through 
    process(BITSEL_u8_u1_7084_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_7084_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_7083_wire_constant = "& Convert_SLV_To_Hex_String(konst_7083_wire_constant) & " outputs:" & " BITSEL_u8_u1_7084_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_7084_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_7084_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7083_wire_constant, tmp_var);
      BITSEL_u8_u1_7084_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_7094_inst flow-through 
    process(BITSEL_u8_u1_7094_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_7094_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_7093_wire_constant = "& Convert_SLV_To_Hex_String(konst_7093_wire_constant) & " outputs:" & " BITSEL_u8_u1_7094_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_7094_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_7094_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7093_wire_constant, tmp_var);
      BITSEL_u8_u1_7094_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_7104_inst flow-through 
    process(BITSEL_u8_u1_7104_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_7104_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_7103_wire_constant = "& Convert_SLV_To_Hex_String(konst_7103_wire_constant) & " outputs:" & " BITSEL_u8_u1_7104_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_7104_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_7104_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7103_wire_constant, tmp_var);
      BITSEL_u8_u1_7104_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_7114_inst flow-through 
    process(BITSEL_u8_u1_7114_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_7114_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_7113_wire_constant = "& Convert_SLV_To_Hex_String(konst_7113_wire_constant) & " outputs:" & " BITSEL_u8_u1_7114_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_7114_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_7114_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7113_wire_constant, tmp_var);
      BITSEL_u8_u1_7114_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_7124_inst flow-through 
    process(BITSEL_u8_u1_7124_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_7124_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_7123_wire_constant = "& Convert_SLV_To_Hex_String(konst_7123_wire_constant) & " outputs:" & " BITSEL_u8_u1_7124_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_7124_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_7124_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7123_wire_constant, tmp_var);
      BITSEL_u8_u1_7124_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_7134_inst flow-through 
    process(BITSEL_u8_u1_7134_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_7134_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_7133_wire_constant = "& Convert_SLV_To_Hex_String(konst_7133_wire_constant) & " outputs:" & " BITSEL_u8_u1_7134_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_7134_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_7134_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7133_wire_constant, tmp_var);
      BITSEL_u8_u1_7134_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_7144_inst flow-through 
    process(BITSEL_u8_u1_7144_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_7144_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_7143_wire_constant = "& Convert_SLV_To_Hex_String(konst_7143_wire_constant) & " outputs:" & " BITSEL_u8_u1_7144_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_7144_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_7144_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7143_wire_constant, tmp_var);
      BITSEL_u8_u1_7144_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_7154_inst flow-through 
    process(BITSEL_u8_u1_7154_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_7154_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_7153_wire_constant = "& Convert_SLV_To_Hex_String(konst_7153_wire_constant) & " outputs:" & " BITSEL_u8_u1_7154_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_7154_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_7154_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7153_wire_constant, tmp_var);
      BITSEL_u8_u1_7154_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_7164_inst flow-through 
    process(BITSEL_u8_u1_7164_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_7164_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_7163_wire_constant = "& Convert_SLV_To_Hex_String(konst_7163_wire_constant) & " outputs:" & " BITSEL_u8_u1_7164_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_7164_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_7164_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7163_wire_constant, tmp_var);
      BITSEL_u8_u1_7164_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_7174_inst flow-through 
    process(BITSEL_u8_u1_7174_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_7174_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_7173_wire_constant = "& Convert_SLV_To_Hex_String(konst_7173_wire_constant) & " outputs:" & " BITSEL_u8_u1_7174_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_7174_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_7174_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7173_wire_constant, tmp_var);
      BITSEL_u8_u1_7174_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_7184_inst flow-through 
    process(BITSEL_u8_u1_7184_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_7184_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_7183_wire_constant = "& Convert_SLV_To_Hex_String(konst_7183_wire_constant) & " outputs:" & " BITSEL_u8_u1_7184_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_7184_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_7184_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7183_wire_constant, tmp_var);
      BITSEL_u8_u1_7184_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_7194_inst flow-through 
    process(BITSEL_u8_u1_7194_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_7194_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_7193_wire_constant = "& Convert_SLV_To_Hex_String(konst_7193_wire_constant) & " outputs:" & " BITSEL_u8_u1_7194_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_7194_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_7194_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7193_wire_constant, tmp_var);
      BITSEL_u8_u1_7194_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_7204_inst flow-through 
    process(BITSEL_u8_u1_7204_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_7204_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_7203_wire_constant = "& Convert_SLV_To_Hex_String(konst_7203_wire_constant) & " outputs:" & " BITSEL_u8_u1_7204_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_7204_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_7204_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7203_wire_constant, tmp_var);
      BITSEL_u8_u1_7204_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_7214_inst flow-through 
    process(BITSEL_u8_u1_7214_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_7214_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_7213_wire_constant = "& Convert_SLV_To_Hex_String(konst_7213_wire_constant) & " outputs:" & " BITSEL_u8_u1_7214_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_7214_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_7214_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7213_wire_constant, tmp_var);
      BITSEL_u8_u1_7214_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_7224_inst flow-through 
    process(BITSEL_u8_u1_7224_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_7224_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_7223_wire_constant = "& Convert_SLV_To_Hex_String(konst_7223_wire_constant) & " outputs:" & " BITSEL_u8_u1_7224_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_7224_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_7224_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7223_wire_constant, tmp_var);
      BITSEL_u8_u1_7224_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_7234_inst flow-through 
    process(BITSEL_u8_u1_7234_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_7234_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_7233_wire_constant = "& Convert_SLV_To_Hex_String(konst_7233_wire_constant) & " outputs:" & " BITSEL_u8_u1_7234_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_7234_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_7234_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7233_wire_constant, tmp_var);
      BITSEL_u8_u1_7234_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_7244_inst flow-through 
    process(BITSEL_u8_u1_7244_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_7244_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_7243_wire_constant = "& Convert_SLV_To_Hex_String(konst_7243_wire_constant) & " outputs:" & " BITSEL_u8_u1_7244_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_7244_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_7244_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7243_wire_constant, tmp_var);
      BITSEL_u8_u1_7244_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_7254_inst flow-through 
    process(BITSEL_u8_u1_7254_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_7254_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_7253_wire_constant = "& Convert_SLV_To_Hex_String(konst_7253_wire_constant) & " outputs:" & " BITSEL_u8_u1_7254_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_7254_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_7254_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7253_wire_constant, tmp_var);
      BITSEL_u8_u1_7254_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_7264_inst flow-through 
    process(BITSEL_u8_u1_7264_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_7264_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_7263_wire_constant = "& Convert_SLV_To_Hex_String(konst_7263_wire_constant) & " outputs:" & " BITSEL_u8_u1_7264_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_7264_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_7264_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7263_wire_constant, tmp_var);
      BITSEL_u8_u1_7264_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_7274_inst flow-through 
    process(BITSEL_u8_u1_7274_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_7274_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_7273_wire_constant = "& Convert_SLV_To_Hex_String(konst_7273_wire_constant) & " outputs:" & " BITSEL_u8_u1_7274_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_7274_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_7274_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7273_wire_constant, tmp_var);
      BITSEL_u8_u1_7274_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_7284_inst flow-through 
    process(BITSEL_u8_u1_7284_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_7284_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_7283_wire_constant = "& Convert_SLV_To_Hex_String(konst_7283_wire_constant) & " outputs:" & " BITSEL_u8_u1_7284_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_7284_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_7284_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7283_wire_constant, tmp_var);
      BITSEL_u8_u1_7284_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_7294_inst flow-through 
    process(BITSEL_u8_u1_7294_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_7294_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_7293_wire_constant = "& Convert_SLV_To_Hex_String(konst_7293_wire_constant) & " outputs:" & " BITSEL_u8_u1_7294_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_7294_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_7294_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7293_wire_constant, tmp_var);
      BITSEL_u8_u1_7294_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_7304_inst flow-through 
    process(BITSEL_u8_u1_7304_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_7304_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_7303_wire_constant = "& Convert_SLV_To_Hex_String(konst_7303_wire_constant) & " outputs:" & " BITSEL_u8_u1_7304_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_7304_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_7304_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7303_wire_constant, tmp_var);
      BITSEL_u8_u1_7304_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_7314_inst flow-through 
    process(BITSEL_u8_u1_7314_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_7314_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_7313_wire_constant = "& Convert_SLV_To_Hex_String(konst_7313_wire_constant) & " outputs:" & " BITSEL_u8_u1_7314_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_7314_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_7314_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7313_wire_constant, tmp_var);
      BITSEL_u8_u1_7314_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_7324_inst flow-through 
    process(BITSEL_u8_u1_7324_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_7324_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_7323_wire_constant = "& Convert_SLV_To_Hex_String(konst_7323_wire_constant) & " outputs:" & " BITSEL_u8_u1_7324_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_7324_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_7324_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7323_wire_constant, tmp_var);
      BITSEL_u8_u1_7324_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_7334_inst flow-through 
    process(BITSEL_u8_u1_7334_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_7334_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_7333_wire_constant = "& Convert_SLV_To_Hex_String(konst_7333_wire_constant) & " outputs:" & " BITSEL_u8_u1_7334_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_7334_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_7334_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7333_wire_constant, tmp_var);
      BITSEL_u8_u1_7334_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_7344_inst flow-through 
    process(BITSEL_u8_u1_7344_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_7344_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_7343_wire_constant = "& Convert_SLV_To_Hex_String(konst_7343_wire_constant) & " outputs:" & " BITSEL_u8_u1_7344_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_7344_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_7344_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7343_wire_constant, tmp_var);
      BITSEL_u8_u1_7344_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_7354_inst flow-through 
    process(BITSEL_u8_u1_7354_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_7354_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_7353_wire_constant = "& Convert_SLV_To_Hex_String(konst_7353_wire_constant) & " outputs:" & " BITSEL_u8_u1_7354_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_7354_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_7354_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7353_wire_constant, tmp_var);
      BITSEL_u8_u1_7354_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_7364_inst flow-through 
    process(BITSEL_u8_u1_7364_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_7364_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_7363_wire_constant = "& Convert_SLV_To_Hex_String(konst_7363_wire_constant) & " outputs:" & " BITSEL_u8_u1_7364_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_7364_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_7364_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7363_wire_constant, tmp_var);
      BITSEL_u8_u1_7364_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_7374_inst flow-through 
    process(BITSEL_u8_u1_7374_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_7374_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_7373_wire_constant = "& Convert_SLV_To_Hex_String(konst_7373_wire_constant) & " outputs:" & " BITSEL_u8_u1_7374_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_7374_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_7374_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7373_wire_constant, tmp_var);
      BITSEL_u8_u1_7374_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_7384_inst flow-through 
    process(BITSEL_u8_u1_7384_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_7384_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_7383_wire_constant = "& Convert_SLV_To_Hex_String(konst_7383_wire_constant) & " outputs:" & " BITSEL_u8_u1_7384_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_7384_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_7384_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7383_wire_constant, tmp_var);
      BITSEL_u8_u1_7384_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_7394_inst flow-through 
    process(BITSEL_u8_u1_7394_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_7394_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_7393_wire_constant = "& Convert_SLV_To_Hex_String(konst_7393_wire_constant) & " outputs:" & " BITSEL_u8_u1_7394_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_7394_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_7394_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7393_wire_constant, tmp_var);
      BITSEL_u8_u1_7394_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_7404_inst flow-through 
    process(BITSEL_u8_u1_7404_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_7404_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_7403_wire_constant = "& Convert_SLV_To_Hex_String(konst_7403_wire_constant) & " outputs:" & " BITSEL_u8_u1_7404_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_7404_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_7404_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7403_wire_constant, tmp_var);
      BITSEL_u8_u1_7404_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_7414_inst flow-through 
    process(BITSEL_u8_u1_7414_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_7414_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_7413_wire_constant = "& Convert_SLV_To_Hex_String(konst_7413_wire_constant) & " outputs:" & " BITSEL_u8_u1_7414_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_7414_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_7414_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7413_wire_constant, tmp_var);
      BITSEL_u8_u1_7414_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_7424_inst flow-through 
    process(BITSEL_u8_u1_7424_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_7424_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_7423_wire_constant = "& Convert_SLV_To_Hex_String(konst_7423_wire_constant) & " outputs:" & " BITSEL_u8_u1_7424_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_7424_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_7424_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7423_wire_constant, tmp_var);
      BITSEL_u8_u1_7424_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_7434_inst flow-through 
    process(BITSEL_u8_u1_7434_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_7434_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_7433_wire_constant = "& Convert_SLV_To_Hex_String(konst_7433_wire_constant) & " outputs:" & " BITSEL_u8_u1_7434_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_7434_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_7434_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7433_wire_constant, tmp_var);
      BITSEL_u8_u1_7434_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_7444_inst flow-through 
    process(BITSEL_u8_u1_7444_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_7444_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_7443_wire_constant = "& Convert_SLV_To_Hex_String(konst_7443_wire_constant) & " outputs:" & " BITSEL_u8_u1_7444_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_7444_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_7444_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7443_wire_constant, tmp_var);
      BITSEL_u8_u1_7444_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_7454_inst flow-through 
    process(BITSEL_u8_u1_7454_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_7454_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_7453_wire_constant = "& Convert_SLV_To_Hex_String(konst_7453_wire_constant) & " outputs:" & " BITSEL_u8_u1_7454_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_7454_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_7454_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7453_wire_constant, tmp_var);
      BITSEL_u8_u1_7454_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_7464_inst flow-through 
    process(BITSEL_u8_u1_7464_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_7464_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_7463_wire_constant = "& Convert_SLV_To_Hex_String(konst_7463_wire_constant) & " outputs:" & " BITSEL_u8_u1_7464_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_7464_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_7464_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7463_wire_constant, tmp_var);
      BITSEL_u8_u1_7464_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_7474_inst flow-through 
    process(BITSEL_u8_u1_7474_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_7474_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_7473_wire_constant = "& Convert_SLV_To_Hex_String(konst_7473_wire_constant) & " outputs:" & " BITSEL_u8_u1_7474_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_7474_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_7474_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7473_wire_constant, tmp_var);
      BITSEL_u8_u1_7474_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_7484_inst flow-through 
    process(BITSEL_u8_u1_7484_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_7484_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_7483_wire_constant = "& Convert_SLV_To_Hex_String(konst_7483_wire_constant) & " outputs:" & " BITSEL_u8_u1_7484_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_7484_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_7484_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7483_wire_constant, tmp_var);
      BITSEL_u8_u1_7484_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_7494_inst flow-through 
    process(BITSEL_u8_u1_7494_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_7494_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_7493_wire_constant = "& Convert_SLV_To_Hex_String(konst_7493_wire_constant) & " outputs:" & " BITSEL_u8_u1_7494_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_7494_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_7494_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7493_wire_constant, tmp_var);
      BITSEL_u8_u1_7494_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_7504_inst flow-through 
    process(BITSEL_u8_u1_7504_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_7504_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_7503_wire_constant = "& Convert_SLV_To_Hex_String(konst_7503_wire_constant) & " outputs:" & " BITSEL_u8_u1_7504_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_7504_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_7504_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7503_wire_constant, tmp_var);
      BITSEL_u8_u1_7504_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_7514_inst flow-through 
    process(BITSEL_u8_u1_7514_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_7514_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_7513_wire_constant = "& Convert_SLV_To_Hex_String(konst_7513_wire_constant) & " outputs:" & " BITSEL_u8_u1_7514_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_7514_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_7514_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7513_wire_constant, tmp_var);
      BITSEL_u8_u1_7514_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_7524_inst flow-through 
    process(BITSEL_u8_u1_7524_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_7524_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_7523_wire_constant = "& Convert_SLV_To_Hex_String(konst_7523_wire_constant) & " outputs:" & " BITSEL_u8_u1_7524_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_7524_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_7524_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7523_wire_constant, tmp_var);
      BITSEL_u8_u1_7524_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_7534_inst flow-through 
    process(BITSEL_u8_u1_7534_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_7534_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_7533_wire_constant = "& Convert_SLV_To_Hex_String(konst_7533_wire_constant) & " outputs:" & " BITSEL_u8_u1_7534_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_7534_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_7534_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7533_wire_constant, tmp_var);
      BITSEL_u8_u1_7534_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_7544_inst flow-through 
    process(BITSEL_u8_u1_7544_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_7544_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_7543_wire_constant = "& Convert_SLV_To_Hex_String(konst_7543_wire_constant) & " outputs:" & " BITSEL_u8_u1_7544_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_7544_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_7544_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7543_wire_constant, tmp_var);
      BITSEL_u8_u1_7544_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_7554_inst flow-through 
    process(BITSEL_u8_u1_7554_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_7554_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_7553_wire_constant = "& Convert_SLV_To_Hex_String(konst_7553_wire_constant) & " outputs:" & " BITSEL_u8_u1_7554_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_7554_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_7554_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7553_wire_constant, tmp_var);
      BITSEL_u8_u1_7554_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_7564_inst flow-through 
    process(BITSEL_u8_u1_7564_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_7564_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_7563_wire_constant = "& Convert_SLV_To_Hex_String(konst_7563_wire_constant) & " outputs:" & " BITSEL_u8_u1_7564_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_7564_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_7564_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7563_wire_constant, tmp_var);
      BITSEL_u8_u1_7564_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_7574_inst flow-through 
    process(BITSEL_u8_u1_7574_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_7574_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_7573_wire_constant = "& Convert_SLV_To_Hex_String(konst_7573_wire_constant) & " outputs:" & " BITSEL_u8_u1_7574_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_7574_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_7574_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7573_wire_constant, tmp_var);
      BITSEL_u8_u1_7574_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_7584_inst flow-through 
    process(BITSEL_u8_u1_7584_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_7584_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_7583_wire_constant = "& Convert_SLV_To_Hex_String(konst_7583_wire_constant) & " outputs:" & " BITSEL_u8_u1_7584_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_7584_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_7584_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7583_wire_constant, tmp_var);
      BITSEL_u8_u1_7584_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_7594_inst flow-through 
    process(BITSEL_u8_u1_7594_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_7594_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_7593_wire_constant = "& Convert_SLV_To_Hex_String(konst_7593_wire_constant) & " outputs:" & " BITSEL_u8_u1_7594_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_7594_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_7594_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7593_wire_constant, tmp_var);
      BITSEL_u8_u1_7594_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_7604_inst flow-through 
    process(BITSEL_u8_u1_7604_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_7604_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_7603_wire_constant = "& Convert_SLV_To_Hex_String(konst_7603_wire_constant) & " outputs:" & " BITSEL_u8_u1_7604_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_7604_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_7604_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7603_wire_constant, tmp_var);
      BITSEL_u8_u1_7604_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_7614_inst flow-through 
    process(BITSEL_u8_u1_7614_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_7614_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_7613_wire_constant = "& Convert_SLV_To_Hex_String(konst_7613_wire_constant) & " outputs:" & " BITSEL_u8_u1_7614_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_7614_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_7614_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7613_wire_constant, tmp_var);
      BITSEL_u8_u1_7614_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_7624_inst flow-through 
    process(BITSEL_u8_u1_7624_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_7624_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_7623_wire_constant = "& Convert_SLV_To_Hex_String(konst_7623_wire_constant) & " outputs:" & " BITSEL_u8_u1_7624_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_7624_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_7624_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7623_wire_constant, tmp_var);
      BITSEL_u8_u1_7624_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_7634_inst flow-through 
    process(BITSEL_u8_u1_7634_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_7634_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_7633_wire_constant = "& Convert_SLV_To_Hex_String(konst_7633_wire_constant) & " outputs:" & " BITSEL_u8_u1_7634_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_7634_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_7634_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7633_wire_constant, tmp_var);
      BITSEL_u8_u1_7634_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_7644_inst flow-through 
    process(BITSEL_u8_u1_7644_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_7644_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_7643_wire_constant = "& Convert_SLV_To_Hex_String(konst_7643_wire_constant) & " outputs:" & " BITSEL_u8_u1_7644_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_7644_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_7644_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7643_wire_constant, tmp_var);
      BITSEL_u8_u1_7644_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_7654_inst flow-through 
    process(BITSEL_u8_u1_7654_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_7654_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_7653_wire_constant = "& Convert_SLV_To_Hex_String(konst_7653_wire_constant) & " outputs:" & " BITSEL_u8_u1_7654_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_7654_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_7654_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7653_wire_constant, tmp_var);
      BITSEL_u8_u1_7654_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_7664_inst flow-through 
    process(BITSEL_u8_u1_7664_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_7664_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_7663_wire_constant = "& Convert_SLV_To_Hex_String(konst_7663_wire_constant) & " outputs:" & " BITSEL_u8_u1_7664_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_7664_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_7664_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7663_wire_constant, tmp_var);
      BITSEL_u8_u1_7664_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_7674_inst flow-through 
    process(BITSEL_u8_u1_7674_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_7674_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_7673_wire_constant = "& Convert_SLV_To_Hex_String(konst_7673_wire_constant) & " outputs:" & " BITSEL_u8_u1_7674_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_7674_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_7674_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7673_wire_constant, tmp_var);
      BITSEL_u8_u1_7674_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_7684_inst flow-through 
    process(BITSEL_u8_u1_7684_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_7684_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_7683_wire_constant = "& Convert_SLV_To_Hex_String(konst_7683_wire_constant) & " outputs:" & " BITSEL_u8_u1_7684_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_7684_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_7684_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7683_wire_constant, tmp_var);
      BITSEL_u8_u1_7684_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_7694_inst flow-through 
    process(BITSEL_u8_u1_7694_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_7694_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_7693_wire_constant = "& Convert_SLV_To_Hex_String(konst_7693_wire_constant) & " outputs:" & " BITSEL_u8_u1_7694_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_7694_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_7694_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7693_wire_constant, tmp_var);
      BITSEL_u8_u1_7694_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_7704_inst flow-through 
    process(BITSEL_u8_u1_7704_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_7704_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_7703_wire_constant = "& Convert_SLV_To_Hex_String(konst_7703_wire_constant) & " outputs:" & " BITSEL_u8_u1_7704_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_7704_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_7704_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7703_wire_constant, tmp_var);
      BITSEL_u8_u1_7704_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_7714_inst flow-through 
    process(BITSEL_u8_u1_7714_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_7714_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_7713_wire_constant = "& Convert_SLV_To_Hex_String(konst_7713_wire_constant) & " outputs:" & " BITSEL_u8_u1_7714_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_7714_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_7714_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7713_wire_constant, tmp_var);
      BITSEL_u8_u1_7714_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_7724_inst flow-through 
    process(BITSEL_u8_u1_7724_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_7724_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_7723_wire_constant = "& Convert_SLV_To_Hex_String(konst_7723_wire_constant) & " outputs:" & " BITSEL_u8_u1_7724_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_7724_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_7724_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7723_wire_constant, tmp_var);
      BITSEL_u8_u1_7724_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_7734_inst flow-through 
    process(BITSEL_u8_u1_7734_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_7734_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_7733_wire_constant = "& Convert_SLV_To_Hex_String(konst_7733_wire_constant) & " outputs:" & " BITSEL_u8_u1_7734_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_7734_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_7734_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7733_wire_constant, tmp_var);
      BITSEL_u8_u1_7734_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_7744_inst flow-through 
    process(BITSEL_u8_u1_7744_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_7744_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_7743_wire_constant = "& Convert_SLV_To_Hex_String(konst_7743_wire_constant) & " outputs:" & " BITSEL_u8_u1_7744_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_7744_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_7744_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7743_wire_constant, tmp_var);
      BITSEL_u8_u1_7744_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_7754_inst flow-through 
    process(BITSEL_u8_u1_7754_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_7754_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_7753_wire_constant = "& Convert_SLV_To_Hex_String(konst_7753_wire_constant) & " outputs:" & " BITSEL_u8_u1_7754_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_7754_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_7754_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7753_wire_constant, tmp_var);
      BITSEL_u8_u1_7754_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_7764_inst flow-through 
    process(BITSEL_u8_u1_7764_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_7764_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_7763_wire_constant = "& Convert_SLV_To_Hex_String(konst_7763_wire_constant) & " outputs:" & " BITSEL_u8_u1_7764_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_7764_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_7764_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7763_wire_constant, tmp_var);
      BITSEL_u8_u1_7764_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_7774_inst flow-through 
    process(BITSEL_u8_u1_7774_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_7774_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_7773_wire_constant = "& Convert_SLV_To_Hex_String(konst_7773_wire_constant) & " outputs:" & " BITSEL_u8_u1_7774_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_7774_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_7774_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7773_wire_constant, tmp_var);
      BITSEL_u8_u1_7774_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_7784_inst flow-through 
    process(BITSEL_u8_u1_7784_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_7784_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_7783_wire_constant = "& Convert_SLV_To_Hex_String(konst_7783_wire_constant) & " outputs:" & " BITSEL_u8_u1_7784_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_7784_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_7784_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7783_wire_constant, tmp_var);
      BITSEL_u8_u1_7784_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_7794_inst flow-through 
    process(BITSEL_u8_u1_7794_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_7794_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_7793_wire_constant = "& Convert_SLV_To_Hex_String(konst_7793_wire_constant) & " outputs:" & " BITSEL_u8_u1_7794_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_7794_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_7794_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7793_wire_constant, tmp_var);
      BITSEL_u8_u1_7794_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_7804_inst flow-through 
    process(BITSEL_u8_u1_7804_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_7804_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_7803_wire_constant = "& Convert_SLV_To_Hex_String(konst_7803_wire_constant) & " outputs:" & " BITSEL_u8_u1_7804_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_7804_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_7804_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7803_wire_constant, tmp_var);
      BITSEL_u8_u1_7804_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_7814_inst flow-through 
    process(BITSEL_u8_u1_7814_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_7814_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_7813_wire_constant = "& Convert_SLV_To_Hex_String(konst_7813_wire_constant) & " outputs:" & " BITSEL_u8_u1_7814_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_7814_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_7814_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7813_wire_constant, tmp_var);
      BITSEL_u8_u1_7814_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_7824_inst flow-through 
    process(BITSEL_u8_u1_7824_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_7824_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_7823_wire_constant = "& Convert_SLV_To_Hex_String(konst_7823_wire_constant) & " outputs:" & " BITSEL_u8_u1_7824_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_7824_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_7824_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7823_wire_constant, tmp_var);
      BITSEL_u8_u1_7824_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_7834_inst flow-through 
    process(BITSEL_u8_u1_7834_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_7834_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_7833_wire_constant = "& Convert_SLV_To_Hex_String(konst_7833_wire_constant) & " outputs:" & " BITSEL_u8_u1_7834_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_7834_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_7834_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7833_wire_constant, tmp_var);
      BITSEL_u8_u1_7834_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_7844_inst flow-through 
    process(BITSEL_u8_u1_7844_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_7844_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_7843_wire_constant = "& Convert_SLV_To_Hex_String(konst_7843_wire_constant) & " outputs:" & " BITSEL_u8_u1_7844_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_7844_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_7844_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7843_wire_constant, tmp_var);
      BITSEL_u8_u1_7844_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_7854_inst flow-through 
    process(BITSEL_u8_u1_7854_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_7854_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_7853_wire_constant = "& Convert_SLV_To_Hex_String(konst_7853_wire_constant) & " outputs:" & " BITSEL_u8_u1_7854_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_7854_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_7854_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7853_wire_constant, tmp_var);
      BITSEL_u8_u1_7854_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_7864_inst flow-through 
    process(BITSEL_u8_u1_7864_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_7864_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_7863_wire_constant = "& Convert_SLV_To_Hex_String(konst_7863_wire_constant) & " outputs:" & " BITSEL_u8_u1_7864_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_7864_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_7864_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7863_wire_constant, tmp_var);
      BITSEL_u8_u1_7864_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_7874_inst flow-through 
    process(BITSEL_u8_u1_7874_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_7874_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_7873_wire_constant = "& Convert_SLV_To_Hex_String(konst_7873_wire_constant) & " outputs:" & " BITSEL_u8_u1_7874_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_7874_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_7874_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7873_wire_constant, tmp_var);
      BITSEL_u8_u1_7874_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_7884_inst flow-through 
    process(BITSEL_u8_u1_7884_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_7884_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_7883_wire_constant = "& Convert_SLV_To_Hex_String(konst_7883_wire_constant) & " outputs:" & " BITSEL_u8_u1_7884_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_7884_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_7884_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7883_wire_constant, tmp_var);
      BITSEL_u8_u1_7884_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_7894_inst flow-through 
    process(BITSEL_u8_u1_7894_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_7894_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_7893_wire_constant = "& Convert_SLV_To_Hex_String(konst_7893_wire_constant) & " outputs:" & " BITSEL_u8_u1_7894_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_7894_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_7894_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7893_wire_constant, tmp_var);
      BITSEL_u8_u1_7894_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_7904_inst flow-through 
    process(BITSEL_u8_u1_7904_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_7904_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_7903_wire_constant = "& Convert_SLV_To_Hex_String(konst_7903_wire_constant) & " outputs:" & " BITSEL_u8_u1_7904_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_7904_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_7904_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7903_wire_constant, tmp_var);
      BITSEL_u8_u1_7904_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_7914_inst flow-through 
    process(BITSEL_u8_u1_7914_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_7914_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_7913_wire_constant = "& Convert_SLV_To_Hex_String(konst_7913_wire_constant) & " outputs:" & " BITSEL_u8_u1_7914_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_7914_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_7914_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7913_wire_constant, tmp_var);
      BITSEL_u8_u1_7914_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_7924_inst flow-through 
    process(BITSEL_u8_u1_7924_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_7924_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_7923_wire_constant = "& Convert_SLV_To_Hex_String(konst_7923_wire_constant) & " outputs:" & " BITSEL_u8_u1_7924_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_7924_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_7924_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7923_wire_constant, tmp_var);
      BITSEL_u8_u1_7924_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_7934_inst flow-through 
    process(BITSEL_u8_u1_7934_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_7934_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_7933_wire_constant = "& Convert_SLV_To_Hex_String(konst_7933_wire_constant) & " outputs:" & " BITSEL_u8_u1_7934_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_7934_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_7934_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7933_wire_constant, tmp_var);
      BITSEL_u8_u1_7934_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_7944_inst flow-through 
    process(BITSEL_u8_u1_7944_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_7944_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_7943_wire_constant = "& Convert_SLV_To_Hex_String(konst_7943_wire_constant) & " outputs:" & " BITSEL_u8_u1_7944_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_7944_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_7944_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7943_wire_constant, tmp_var);
      BITSEL_u8_u1_7944_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_7954_inst flow-through 
    process(BITSEL_u8_u1_7954_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_7954_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_7953_wire_constant = "& Convert_SLV_To_Hex_String(konst_7953_wire_constant) & " outputs:" & " BITSEL_u8_u1_7954_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_7954_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_7954_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7953_wire_constant, tmp_var);
      BITSEL_u8_u1_7954_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_7964_inst flow-through 
    process(BITSEL_u8_u1_7964_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_7964_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_7963_wire_constant = "& Convert_SLV_To_Hex_String(konst_7963_wire_constant) & " outputs:" & " BITSEL_u8_u1_7964_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_7964_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_7964_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7963_wire_constant, tmp_var);
      BITSEL_u8_u1_7964_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_7974_inst flow-through 
    process(BITSEL_u8_u1_7974_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_7974_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_7973_wire_constant = "& Convert_SLV_To_Hex_String(konst_7973_wire_constant) & " outputs:" & " BITSEL_u8_u1_7974_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_7974_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_7974_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7973_wire_constant, tmp_var);
      BITSEL_u8_u1_7974_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_7984_inst flow-through 
    process(BITSEL_u8_u1_7984_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_7984_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_7983_wire_constant = "& Convert_SLV_To_Hex_String(konst_7983_wire_constant) & " outputs:" & " BITSEL_u8_u1_7984_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_7984_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_7984_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7983_wire_constant, tmp_var);
      BITSEL_u8_u1_7984_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_7994_inst flow-through 
    process(BITSEL_u8_u1_7994_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_7994_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_7993_wire_constant = "& Convert_SLV_To_Hex_String(konst_7993_wire_constant) & " outputs:" & " BITSEL_u8_u1_7994_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_7994_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_7994_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7993_wire_constant, tmp_var);
      BITSEL_u8_u1_7994_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8004_inst flow-through 
    process(BITSEL_u8_u1_8004_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8004_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8003_wire_constant = "& Convert_SLV_To_Hex_String(konst_8003_wire_constant) & " outputs:" & " BITSEL_u8_u1_8004_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8004_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8004_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8003_wire_constant, tmp_var);
      BITSEL_u8_u1_8004_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8014_inst flow-through 
    process(BITSEL_u8_u1_8014_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8014_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8013_wire_constant = "& Convert_SLV_To_Hex_String(konst_8013_wire_constant) & " outputs:" & " BITSEL_u8_u1_8014_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8014_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8014_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8013_wire_constant, tmp_var);
      BITSEL_u8_u1_8014_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8024_inst flow-through 
    process(BITSEL_u8_u1_8024_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8024_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8023_wire_constant = "& Convert_SLV_To_Hex_String(konst_8023_wire_constant) & " outputs:" & " BITSEL_u8_u1_8024_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8024_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8024_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8023_wire_constant, tmp_var);
      BITSEL_u8_u1_8024_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8034_inst flow-through 
    process(BITSEL_u8_u1_8034_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8034_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8033_wire_constant = "& Convert_SLV_To_Hex_String(konst_8033_wire_constant) & " outputs:" & " BITSEL_u8_u1_8034_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8034_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8034_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8033_wire_constant, tmp_var);
      BITSEL_u8_u1_8034_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8044_inst flow-through 
    process(BITSEL_u8_u1_8044_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8044_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8043_wire_constant = "& Convert_SLV_To_Hex_String(konst_8043_wire_constant) & " outputs:" & " BITSEL_u8_u1_8044_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8044_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8044_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8043_wire_constant, tmp_var);
      BITSEL_u8_u1_8044_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8054_inst flow-through 
    process(BITSEL_u8_u1_8054_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8054_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8053_wire_constant = "& Convert_SLV_To_Hex_String(konst_8053_wire_constant) & " outputs:" & " BITSEL_u8_u1_8054_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8054_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8054_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8053_wire_constant, tmp_var);
      BITSEL_u8_u1_8054_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8064_inst flow-through 
    process(BITSEL_u8_u1_8064_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8064_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8063_wire_constant = "& Convert_SLV_To_Hex_String(konst_8063_wire_constant) & " outputs:" & " BITSEL_u8_u1_8064_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8064_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8064_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8063_wire_constant, tmp_var);
      BITSEL_u8_u1_8064_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8074_inst flow-through 
    process(BITSEL_u8_u1_8074_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8074_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8073_wire_constant = "& Convert_SLV_To_Hex_String(konst_8073_wire_constant) & " outputs:" & " BITSEL_u8_u1_8074_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8074_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8074_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8073_wire_constant, tmp_var);
      BITSEL_u8_u1_8074_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8084_inst flow-through 
    process(BITSEL_u8_u1_8084_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8084_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8083_wire_constant = "& Convert_SLV_To_Hex_String(konst_8083_wire_constant) & " outputs:" & " BITSEL_u8_u1_8084_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8084_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8084_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8083_wire_constant, tmp_var);
      BITSEL_u8_u1_8084_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8094_inst flow-through 
    process(BITSEL_u8_u1_8094_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8094_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8093_wire_constant = "& Convert_SLV_To_Hex_String(konst_8093_wire_constant) & " outputs:" & " BITSEL_u8_u1_8094_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8094_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8094_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8093_wire_constant, tmp_var);
      BITSEL_u8_u1_8094_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8104_inst flow-through 
    process(BITSEL_u8_u1_8104_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8104_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8103_wire_constant = "& Convert_SLV_To_Hex_String(konst_8103_wire_constant) & " outputs:" & " BITSEL_u8_u1_8104_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8104_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8104_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8103_wire_constant, tmp_var);
      BITSEL_u8_u1_8104_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8114_inst flow-through 
    process(BITSEL_u8_u1_8114_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8114_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8113_wire_constant = "& Convert_SLV_To_Hex_String(konst_8113_wire_constant) & " outputs:" & " BITSEL_u8_u1_8114_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8114_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8114_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8113_wire_constant, tmp_var);
      BITSEL_u8_u1_8114_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8124_inst flow-through 
    process(BITSEL_u8_u1_8124_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8124_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8123_wire_constant = "& Convert_SLV_To_Hex_String(konst_8123_wire_constant) & " outputs:" & " BITSEL_u8_u1_8124_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8124_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8124_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8123_wire_constant, tmp_var);
      BITSEL_u8_u1_8124_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8134_inst flow-through 
    process(BITSEL_u8_u1_8134_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8134_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8133_wire_constant = "& Convert_SLV_To_Hex_String(konst_8133_wire_constant) & " outputs:" & " BITSEL_u8_u1_8134_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8134_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8134_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8133_wire_constant, tmp_var);
      BITSEL_u8_u1_8134_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8144_inst flow-through 
    process(BITSEL_u8_u1_8144_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8144_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8143_wire_constant = "& Convert_SLV_To_Hex_String(konst_8143_wire_constant) & " outputs:" & " BITSEL_u8_u1_8144_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8144_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8144_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8143_wire_constant, tmp_var);
      BITSEL_u8_u1_8144_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8154_inst flow-through 
    process(BITSEL_u8_u1_8154_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8154_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8153_wire_constant = "& Convert_SLV_To_Hex_String(konst_8153_wire_constant) & " outputs:" & " BITSEL_u8_u1_8154_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8154_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8154_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8153_wire_constant, tmp_var);
      BITSEL_u8_u1_8154_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8164_inst flow-through 
    process(BITSEL_u8_u1_8164_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8164_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8163_wire_constant = "& Convert_SLV_To_Hex_String(konst_8163_wire_constant) & " outputs:" & " BITSEL_u8_u1_8164_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8164_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8164_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8163_wire_constant, tmp_var);
      BITSEL_u8_u1_8164_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8174_inst flow-through 
    process(BITSEL_u8_u1_8174_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8174_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8173_wire_constant = "& Convert_SLV_To_Hex_String(konst_8173_wire_constant) & " outputs:" & " BITSEL_u8_u1_8174_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8174_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8174_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8173_wire_constant, tmp_var);
      BITSEL_u8_u1_8174_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8184_inst flow-through 
    process(BITSEL_u8_u1_8184_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8184_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8183_wire_constant = "& Convert_SLV_To_Hex_String(konst_8183_wire_constant) & " outputs:" & " BITSEL_u8_u1_8184_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8184_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8184_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8183_wire_constant, tmp_var);
      BITSEL_u8_u1_8184_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8194_inst flow-through 
    process(BITSEL_u8_u1_8194_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8194_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8193_wire_constant = "& Convert_SLV_To_Hex_String(konst_8193_wire_constant) & " outputs:" & " BITSEL_u8_u1_8194_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8194_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8194_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8193_wire_constant, tmp_var);
      BITSEL_u8_u1_8194_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8202_inst flow-through 
    process(BITSEL_u8_u1_8202_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8202_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8201_wire_constant = "& Convert_SLV_To_Hex_String(konst_8201_wire_constant) & " outputs:" & " BITSEL_u8_u1_8202_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8202_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8202_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8201_wire_constant, tmp_var);
      BITSEL_u8_u1_8202_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8210_inst flow-through 
    process(BITSEL_u8_u1_8210_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8210_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8209_wire_constant = "& Convert_SLV_To_Hex_String(konst_8209_wire_constant) & " outputs:" & " BITSEL_u8_u1_8210_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8210_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8210_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8209_wire_constant, tmp_var);
      BITSEL_u8_u1_8210_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8218_inst flow-through 
    process(BITSEL_u8_u1_8218_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8218_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8217_wire_constant = "& Convert_SLV_To_Hex_String(konst_8217_wire_constant) & " outputs:" & " BITSEL_u8_u1_8218_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8218_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8218_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8217_wire_constant, tmp_var);
      BITSEL_u8_u1_8218_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8226_inst flow-through 
    process(BITSEL_u8_u1_8226_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8226_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8225_wire_constant = "& Convert_SLV_To_Hex_String(konst_8225_wire_constant) & " outputs:" & " BITSEL_u8_u1_8226_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8226_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8226_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8225_wire_constant, tmp_var);
      BITSEL_u8_u1_8226_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8234_inst flow-through 
    process(BITSEL_u8_u1_8234_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8234_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8233_wire_constant = "& Convert_SLV_To_Hex_String(konst_8233_wire_constant) & " outputs:" & " BITSEL_u8_u1_8234_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8234_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8234_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8233_wire_constant, tmp_var);
      BITSEL_u8_u1_8234_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8242_inst flow-through 
    process(BITSEL_u8_u1_8242_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8242_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8241_wire_constant = "& Convert_SLV_To_Hex_String(konst_8241_wire_constant) & " outputs:" & " BITSEL_u8_u1_8242_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8242_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8242_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8241_wire_constant, tmp_var);
      BITSEL_u8_u1_8242_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8250_inst flow-through 
    process(BITSEL_u8_u1_8250_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8250_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8249_wire_constant = "& Convert_SLV_To_Hex_String(konst_8249_wire_constant) & " outputs:" & " BITSEL_u8_u1_8250_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8250_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8250_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8249_wire_constant, tmp_var);
      BITSEL_u8_u1_8250_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8258_inst flow-through 
    process(BITSEL_u8_u1_8258_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8258_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8257_wire_constant = "& Convert_SLV_To_Hex_String(konst_8257_wire_constant) & " outputs:" & " BITSEL_u8_u1_8258_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8258_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8258_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8257_wire_constant, tmp_var);
      BITSEL_u8_u1_8258_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8266_inst flow-through 
    process(BITSEL_u8_u1_8266_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8266_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8265_wire_constant = "& Convert_SLV_To_Hex_String(konst_8265_wire_constant) & " outputs:" & " BITSEL_u8_u1_8266_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8266_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8266_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8265_wire_constant, tmp_var);
      BITSEL_u8_u1_8266_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8274_inst flow-through 
    process(BITSEL_u8_u1_8274_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8274_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8273_wire_constant = "& Convert_SLV_To_Hex_String(konst_8273_wire_constant) & " outputs:" & " BITSEL_u8_u1_8274_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8274_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8274_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8273_wire_constant, tmp_var);
      BITSEL_u8_u1_8274_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8282_inst flow-through 
    process(BITSEL_u8_u1_8282_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8282_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8281_wire_constant = "& Convert_SLV_To_Hex_String(konst_8281_wire_constant) & " outputs:" & " BITSEL_u8_u1_8282_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8282_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8282_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8281_wire_constant, tmp_var);
      BITSEL_u8_u1_8282_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8290_inst flow-through 
    process(BITSEL_u8_u1_8290_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8290_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8289_wire_constant = "& Convert_SLV_To_Hex_String(konst_8289_wire_constant) & " outputs:" & " BITSEL_u8_u1_8290_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8290_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8290_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8289_wire_constant, tmp_var);
      BITSEL_u8_u1_8290_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8298_inst flow-through 
    process(BITSEL_u8_u1_8298_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8298_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8297_wire_constant = "& Convert_SLV_To_Hex_String(konst_8297_wire_constant) & " outputs:" & " BITSEL_u8_u1_8298_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8298_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8298_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8297_wire_constant, tmp_var);
      BITSEL_u8_u1_8298_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8306_inst flow-through 
    process(BITSEL_u8_u1_8306_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8306_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8305_wire_constant = "& Convert_SLV_To_Hex_String(konst_8305_wire_constant) & " outputs:" & " BITSEL_u8_u1_8306_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8306_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8306_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8305_wire_constant, tmp_var);
      BITSEL_u8_u1_8306_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8314_inst flow-through 
    process(BITSEL_u8_u1_8314_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8314_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8313_wire_constant = "& Convert_SLV_To_Hex_String(konst_8313_wire_constant) & " outputs:" & " BITSEL_u8_u1_8314_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8314_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8314_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8313_wire_constant, tmp_var);
      BITSEL_u8_u1_8314_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8322_inst flow-through 
    process(BITSEL_u8_u1_8322_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8322_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8321_wire_constant = "& Convert_SLV_To_Hex_String(konst_8321_wire_constant) & " outputs:" & " BITSEL_u8_u1_8322_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8322_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8322_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8321_wire_constant, tmp_var);
      BITSEL_u8_u1_8322_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8330_inst flow-through 
    process(BITSEL_u8_u1_8330_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8330_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8329_wire_constant = "& Convert_SLV_To_Hex_String(konst_8329_wire_constant) & " outputs:" & " BITSEL_u8_u1_8330_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8330_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8330_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8329_wire_constant, tmp_var);
      BITSEL_u8_u1_8330_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8338_inst flow-through 
    process(BITSEL_u8_u1_8338_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8338_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8337_wire_constant = "& Convert_SLV_To_Hex_String(konst_8337_wire_constant) & " outputs:" & " BITSEL_u8_u1_8338_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8338_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8338_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8337_wire_constant, tmp_var);
      BITSEL_u8_u1_8338_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8346_inst flow-through 
    process(BITSEL_u8_u1_8346_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8346_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8345_wire_constant = "& Convert_SLV_To_Hex_String(konst_8345_wire_constant) & " outputs:" & " BITSEL_u8_u1_8346_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8346_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8346_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8345_wire_constant, tmp_var);
      BITSEL_u8_u1_8346_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8354_inst flow-through 
    process(BITSEL_u8_u1_8354_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8354_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8353_wire_constant = "& Convert_SLV_To_Hex_String(konst_8353_wire_constant) & " outputs:" & " BITSEL_u8_u1_8354_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8354_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8354_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8353_wire_constant, tmp_var);
      BITSEL_u8_u1_8354_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8362_inst flow-through 
    process(BITSEL_u8_u1_8362_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8362_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8361_wire_constant = "& Convert_SLV_To_Hex_String(konst_8361_wire_constant) & " outputs:" & " BITSEL_u8_u1_8362_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8362_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8362_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8361_wire_constant, tmp_var);
      BITSEL_u8_u1_8362_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8370_inst flow-through 
    process(BITSEL_u8_u1_8370_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8370_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8369_wire_constant = "& Convert_SLV_To_Hex_String(konst_8369_wire_constant) & " outputs:" & " BITSEL_u8_u1_8370_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8370_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8370_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8369_wire_constant, tmp_var);
      BITSEL_u8_u1_8370_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8378_inst flow-through 
    process(BITSEL_u8_u1_8378_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8378_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8377_wire_constant = "& Convert_SLV_To_Hex_String(konst_8377_wire_constant) & " outputs:" & " BITSEL_u8_u1_8378_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8378_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8378_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8377_wire_constant, tmp_var);
      BITSEL_u8_u1_8378_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8386_inst flow-through 
    process(BITSEL_u8_u1_8386_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8386_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8385_wire_constant = "& Convert_SLV_To_Hex_String(konst_8385_wire_constant) & " outputs:" & " BITSEL_u8_u1_8386_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8386_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8386_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8385_wire_constant, tmp_var);
      BITSEL_u8_u1_8386_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8394_inst flow-through 
    process(BITSEL_u8_u1_8394_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8394_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8393_wire_constant = "& Convert_SLV_To_Hex_String(konst_8393_wire_constant) & " outputs:" & " BITSEL_u8_u1_8394_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8394_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8394_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8393_wire_constant, tmp_var);
      BITSEL_u8_u1_8394_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8402_inst flow-through 
    process(BITSEL_u8_u1_8402_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8402_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8401_wire_constant = "& Convert_SLV_To_Hex_String(konst_8401_wire_constant) & " outputs:" & " BITSEL_u8_u1_8402_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8402_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8402_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8401_wire_constant, tmp_var);
      BITSEL_u8_u1_8402_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8410_inst flow-through 
    process(BITSEL_u8_u1_8410_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8410_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8409_wire_constant = "& Convert_SLV_To_Hex_String(konst_8409_wire_constant) & " outputs:" & " BITSEL_u8_u1_8410_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8410_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8410_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8409_wire_constant, tmp_var);
      BITSEL_u8_u1_8410_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8418_inst flow-through 
    process(BITSEL_u8_u1_8418_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8418_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8417_wire_constant = "& Convert_SLV_To_Hex_String(konst_8417_wire_constant) & " outputs:" & " BITSEL_u8_u1_8418_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8418_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8418_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8417_wire_constant, tmp_var);
      BITSEL_u8_u1_8418_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8426_inst flow-through 
    process(BITSEL_u8_u1_8426_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8426_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8425_wire_constant = "& Convert_SLV_To_Hex_String(konst_8425_wire_constant) & " outputs:" & " BITSEL_u8_u1_8426_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8426_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8426_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8425_wire_constant, tmp_var);
      BITSEL_u8_u1_8426_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8434_inst flow-through 
    process(BITSEL_u8_u1_8434_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8434_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8433_wire_constant = "& Convert_SLV_To_Hex_String(konst_8433_wire_constant) & " outputs:" & " BITSEL_u8_u1_8434_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8434_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8434_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8433_wire_constant, tmp_var);
      BITSEL_u8_u1_8434_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8442_inst flow-through 
    process(BITSEL_u8_u1_8442_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8442_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8441_wire_constant = "& Convert_SLV_To_Hex_String(konst_8441_wire_constant) & " outputs:" & " BITSEL_u8_u1_8442_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8442_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8442_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8441_wire_constant, tmp_var);
      BITSEL_u8_u1_8442_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8450_inst flow-through 
    process(BITSEL_u8_u1_8450_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8450_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8449_wire_constant = "& Convert_SLV_To_Hex_String(konst_8449_wire_constant) & " outputs:" & " BITSEL_u8_u1_8450_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8450_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8450_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8449_wire_constant, tmp_var);
      BITSEL_u8_u1_8450_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8458_inst flow-through 
    process(BITSEL_u8_u1_8458_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8458_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8457_wire_constant = "& Convert_SLV_To_Hex_String(konst_8457_wire_constant) & " outputs:" & " BITSEL_u8_u1_8458_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8458_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8458_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8457_wire_constant, tmp_var);
      BITSEL_u8_u1_8458_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8466_inst flow-through 
    process(BITSEL_u8_u1_8466_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8466_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8465_wire_constant = "& Convert_SLV_To_Hex_String(konst_8465_wire_constant) & " outputs:" & " BITSEL_u8_u1_8466_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8466_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8466_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8465_wire_constant, tmp_var);
      BITSEL_u8_u1_8466_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8474_inst flow-through 
    process(BITSEL_u8_u1_8474_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8474_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8473_wire_constant = "& Convert_SLV_To_Hex_String(konst_8473_wire_constant) & " outputs:" & " BITSEL_u8_u1_8474_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8474_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8474_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8473_wire_constant, tmp_var);
      BITSEL_u8_u1_8474_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8482_inst flow-through 
    process(BITSEL_u8_u1_8482_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8482_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8481_wire_constant = "& Convert_SLV_To_Hex_String(konst_8481_wire_constant) & " outputs:" & " BITSEL_u8_u1_8482_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8482_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8482_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8481_wire_constant, tmp_var);
      BITSEL_u8_u1_8482_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8490_inst flow-through 
    process(BITSEL_u8_u1_8490_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8490_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8489_wire_constant = "& Convert_SLV_To_Hex_String(konst_8489_wire_constant) & " outputs:" & " BITSEL_u8_u1_8490_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8490_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8490_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8489_wire_constant, tmp_var);
      BITSEL_u8_u1_8490_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8498_inst flow-through 
    process(BITSEL_u8_u1_8498_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8498_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8497_wire_constant = "& Convert_SLV_To_Hex_String(konst_8497_wire_constant) & " outputs:" & " BITSEL_u8_u1_8498_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8498_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8498_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8497_wire_constant, tmp_var);
      BITSEL_u8_u1_8498_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8506_inst flow-through 
    process(BITSEL_u8_u1_8506_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8506_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8505_wire_constant = "& Convert_SLV_To_Hex_String(konst_8505_wire_constant) & " outputs:" & " BITSEL_u8_u1_8506_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8506_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8506_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8505_wire_constant, tmp_var);
      BITSEL_u8_u1_8506_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8514_inst flow-through 
    process(BITSEL_u8_u1_8514_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8514_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8513_wire_constant = "& Convert_SLV_To_Hex_String(konst_8513_wire_constant) & " outputs:" & " BITSEL_u8_u1_8514_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8514_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8514_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8513_wire_constant, tmp_var);
      BITSEL_u8_u1_8514_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8522_inst flow-through 
    process(BITSEL_u8_u1_8522_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8522_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8521_wire_constant = "& Convert_SLV_To_Hex_String(konst_8521_wire_constant) & " outputs:" & " BITSEL_u8_u1_8522_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8522_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8522_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8521_wire_constant, tmp_var);
      BITSEL_u8_u1_8522_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8530_inst flow-through 
    process(BITSEL_u8_u1_8530_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8530_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8529_wire_constant = "& Convert_SLV_To_Hex_String(konst_8529_wire_constant) & " outputs:" & " BITSEL_u8_u1_8530_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8530_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8530_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8529_wire_constant, tmp_var);
      BITSEL_u8_u1_8530_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8538_inst flow-through 
    process(BITSEL_u8_u1_8538_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8538_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8537_wire_constant = "& Convert_SLV_To_Hex_String(konst_8537_wire_constant) & " outputs:" & " BITSEL_u8_u1_8538_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8538_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8538_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8537_wire_constant, tmp_var);
      BITSEL_u8_u1_8538_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8546_inst flow-through 
    process(BITSEL_u8_u1_8546_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8546_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8545_wire_constant = "& Convert_SLV_To_Hex_String(konst_8545_wire_constant) & " outputs:" & " BITSEL_u8_u1_8546_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8546_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8546_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8545_wire_constant, tmp_var);
      BITSEL_u8_u1_8546_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8554_inst flow-through 
    process(BITSEL_u8_u1_8554_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8554_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8553_wire_constant = "& Convert_SLV_To_Hex_String(konst_8553_wire_constant) & " outputs:" & " BITSEL_u8_u1_8554_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8554_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8554_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8553_wire_constant, tmp_var);
      BITSEL_u8_u1_8554_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8562_inst flow-through 
    process(BITSEL_u8_u1_8562_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8562_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8561_wire_constant = "& Convert_SLV_To_Hex_String(konst_8561_wire_constant) & " outputs:" & " BITSEL_u8_u1_8562_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8562_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8562_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8561_wire_constant, tmp_var);
      BITSEL_u8_u1_8562_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8570_inst flow-through 
    process(BITSEL_u8_u1_8570_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8570_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8569_wire_constant = "& Convert_SLV_To_Hex_String(konst_8569_wire_constant) & " outputs:" & " BITSEL_u8_u1_8570_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8570_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8570_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8569_wire_constant, tmp_var);
      BITSEL_u8_u1_8570_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8578_inst flow-through 
    process(BITSEL_u8_u1_8578_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8578_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8577_wire_constant = "& Convert_SLV_To_Hex_String(konst_8577_wire_constant) & " outputs:" & " BITSEL_u8_u1_8578_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8578_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8578_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8577_wire_constant, tmp_var);
      BITSEL_u8_u1_8578_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8586_inst flow-through 
    process(BITSEL_u8_u1_8586_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8586_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8585_wire_constant = "& Convert_SLV_To_Hex_String(konst_8585_wire_constant) & " outputs:" & " BITSEL_u8_u1_8586_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8586_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8586_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8585_wire_constant, tmp_var);
      BITSEL_u8_u1_8586_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8594_inst flow-through 
    process(BITSEL_u8_u1_8594_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8594_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8593_wire_constant = "& Convert_SLV_To_Hex_String(konst_8593_wire_constant) & " outputs:" & " BITSEL_u8_u1_8594_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8594_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8594_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8593_wire_constant, tmp_var);
      BITSEL_u8_u1_8594_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8602_inst flow-through 
    process(BITSEL_u8_u1_8602_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8602_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8601_wire_constant = "& Convert_SLV_To_Hex_String(konst_8601_wire_constant) & " outputs:" & " BITSEL_u8_u1_8602_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8602_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8602_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8601_wire_constant, tmp_var);
      BITSEL_u8_u1_8602_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8610_inst flow-through 
    process(BITSEL_u8_u1_8610_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8610_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8609_wire_constant = "& Convert_SLV_To_Hex_String(konst_8609_wire_constant) & " outputs:" & " BITSEL_u8_u1_8610_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8610_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8610_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8609_wire_constant, tmp_var);
      BITSEL_u8_u1_8610_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8618_inst flow-through 
    process(BITSEL_u8_u1_8618_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8618_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8617_wire_constant = "& Convert_SLV_To_Hex_String(konst_8617_wire_constant) & " outputs:" & " BITSEL_u8_u1_8618_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8618_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8618_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8617_wire_constant, tmp_var);
      BITSEL_u8_u1_8618_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8626_inst flow-through 
    process(BITSEL_u8_u1_8626_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8626_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8625_wire_constant = "& Convert_SLV_To_Hex_String(konst_8625_wire_constant) & " outputs:" & " BITSEL_u8_u1_8626_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8626_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8626_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8625_wire_constant, tmp_var);
      BITSEL_u8_u1_8626_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8634_inst flow-through 
    process(BITSEL_u8_u1_8634_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8634_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8633_wire_constant = "& Convert_SLV_To_Hex_String(konst_8633_wire_constant) & " outputs:" & " BITSEL_u8_u1_8634_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8634_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8634_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8633_wire_constant, tmp_var);
      BITSEL_u8_u1_8634_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8642_inst flow-through 
    process(BITSEL_u8_u1_8642_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8642_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8641_wire_constant = "& Convert_SLV_To_Hex_String(konst_8641_wire_constant) & " outputs:" & " BITSEL_u8_u1_8642_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8642_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8642_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8641_wire_constant, tmp_var);
      BITSEL_u8_u1_8642_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8650_inst flow-through 
    process(BITSEL_u8_u1_8650_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8650_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8649_wire_constant = "& Convert_SLV_To_Hex_String(konst_8649_wire_constant) & " outputs:" & " BITSEL_u8_u1_8650_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8650_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8650_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8649_wire_constant, tmp_var);
      BITSEL_u8_u1_8650_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8658_inst flow-through 
    process(BITSEL_u8_u1_8658_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8658_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8657_wire_constant = "& Convert_SLV_To_Hex_String(konst_8657_wire_constant) & " outputs:" & " BITSEL_u8_u1_8658_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8658_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8658_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8657_wire_constant, tmp_var);
      BITSEL_u8_u1_8658_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8666_inst flow-through 
    process(BITSEL_u8_u1_8666_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8666_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8665_wire_constant = "& Convert_SLV_To_Hex_String(konst_8665_wire_constant) & " outputs:" & " BITSEL_u8_u1_8666_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8666_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8666_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8665_wire_constant, tmp_var);
      BITSEL_u8_u1_8666_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8674_inst flow-through 
    process(BITSEL_u8_u1_8674_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8674_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8673_wire_constant = "& Convert_SLV_To_Hex_String(konst_8673_wire_constant) & " outputs:" & " BITSEL_u8_u1_8674_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8674_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8674_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8673_wire_constant, tmp_var);
      BITSEL_u8_u1_8674_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8682_inst flow-through 
    process(BITSEL_u8_u1_8682_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8682_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8681_wire_constant = "& Convert_SLV_To_Hex_String(konst_8681_wire_constant) & " outputs:" & " BITSEL_u8_u1_8682_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8682_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8682_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8681_wire_constant, tmp_var);
      BITSEL_u8_u1_8682_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8690_inst flow-through 
    process(BITSEL_u8_u1_8690_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8690_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8689_wire_constant = "& Convert_SLV_To_Hex_String(konst_8689_wire_constant) & " outputs:" & " BITSEL_u8_u1_8690_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8690_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8690_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8689_wire_constant, tmp_var);
      BITSEL_u8_u1_8690_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8698_inst flow-through 
    process(BITSEL_u8_u1_8698_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8698_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8697_wire_constant = "& Convert_SLV_To_Hex_String(konst_8697_wire_constant) & " outputs:" & " BITSEL_u8_u1_8698_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8698_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8698_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8697_wire_constant, tmp_var);
      BITSEL_u8_u1_8698_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8706_inst flow-through 
    process(BITSEL_u8_u1_8706_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8706_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8705_wire_constant = "& Convert_SLV_To_Hex_String(konst_8705_wire_constant) & " outputs:" & " BITSEL_u8_u1_8706_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8706_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8706_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8705_wire_constant, tmp_var);
      BITSEL_u8_u1_8706_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8714_inst flow-through 
    process(BITSEL_u8_u1_8714_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8714_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8713_wire_constant = "& Convert_SLV_To_Hex_String(konst_8713_wire_constant) & " outputs:" & " BITSEL_u8_u1_8714_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8714_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8714_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8713_wire_constant, tmp_var);
      BITSEL_u8_u1_8714_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8722_inst flow-through 
    process(BITSEL_u8_u1_8722_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8722_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8721_wire_constant = "& Convert_SLV_To_Hex_String(konst_8721_wire_constant) & " outputs:" & " BITSEL_u8_u1_8722_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8722_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8722_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8721_wire_constant, tmp_var);
      BITSEL_u8_u1_8722_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8730_inst flow-through 
    process(BITSEL_u8_u1_8730_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8730_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8729_wire_constant = "& Convert_SLV_To_Hex_String(konst_8729_wire_constant) & " outputs:" & " BITSEL_u8_u1_8730_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8730_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8730_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8729_wire_constant, tmp_var);
      BITSEL_u8_u1_8730_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8738_inst flow-through 
    process(BITSEL_u8_u1_8738_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8738_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8737_wire_constant = "& Convert_SLV_To_Hex_String(konst_8737_wire_constant) & " outputs:" & " BITSEL_u8_u1_8738_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8738_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8738_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8737_wire_constant, tmp_var);
      BITSEL_u8_u1_8738_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8746_inst flow-through 
    process(BITSEL_u8_u1_8746_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8746_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8745_wire_constant = "& Convert_SLV_To_Hex_String(konst_8745_wire_constant) & " outputs:" & " BITSEL_u8_u1_8746_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8746_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8746_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8745_wire_constant, tmp_var);
      BITSEL_u8_u1_8746_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8754_inst flow-through 
    process(BITSEL_u8_u1_8754_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8754_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8753_wire_constant = "& Convert_SLV_To_Hex_String(konst_8753_wire_constant) & " outputs:" & " BITSEL_u8_u1_8754_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8754_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8754_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8753_wire_constant, tmp_var);
      BITSEL_u8_u1_8754_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8762_inst flow-through 
    process(BITSEL_u8_u1_8762_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8762_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8761_wire_constant = "& Convert_SLV_To_Hex_String(konst_8761_wire_constant) & " outputs:" & " BITSEL_u8_u1_8762_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8762_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8762_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8761_wire_constant, tmp_var);
      BITSEL_u8_u1_8762_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8770_inst flow-through 
    process(BITSEL_u8_u1_8770_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8770_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8769_wire_constant = "& Convert_SLV_To_Hex_String(konst_8769_wire_constant) & " outputs:" & " BITSEL_u8_u1_8770_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8770_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8770_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8769_wire_constant, tmp_var);
      BITSEL_u8_u1_8770_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8778_inst flow-through 
    process(BITSEL_u8_u1_8778_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8778_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8777_wire_constant = "& Convert_SLV_To_Hex_String(konst_8777_wire_constant) & " outputs:" & " BITSEL_u8_u1_8778_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8778_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8778_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8777_wire_constant, tmp_var);
      BITSEL_u8_u1_8778_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8786_inst flow-through 
    process(BITSEL_u8_u1_8786_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8786_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8785_wire_constant = "& Convert_SLV_To_Hex_String(konst_8785_wire_constant) & " outputs:" & " BITSEL_u8_u1_8786_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8786_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8786_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8785_wire_constant, tmp_var);
      BITSEL_u8_u1_8786_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8794_inst flow-through 
    process(BITSEL_u8_u1_8794_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8794_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8793_wire_constant = "& Convert_SLV_To_Hex_String(konst_8793_wire_constant) & " outputs:" & " BITSEL_u8_u1_8794_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8794_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8794_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8793_wire_constant, tmp_var);
      BITSEL_u8_u1_8794_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8802_inst flow-through 
    process(BITSEL_u8_u1_8802_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8802_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8801_wire_constant = "& Convert_SLV_To_Hex_String(konst_8801_wire_constant) & " outputs:" & " BITSEL_u8_u1_8802_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8802_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8802_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8801_wire_constant, tmp_var);
      BITSEL_u8_u1_8802_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8810_inst flow-through 
    process(BITSEL_u8_u1_8810_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8810_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8809_wire_constant = "& Convert_SLV_To_Hex_String(konst_8809_wire_constant) & " outputs:" & " BITSEL_u8_u1_8810_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8810_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8810_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8809_wire_constant, tmp_var);
      BITSEL_u8_u1_8810_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8818_inst flow-through 
    process(BITSEL_u8_u1_8818_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8818_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8817_wire_constant = "& Convert_SLV_To_Hex_String(konst_8817_wire_constant) & " outputs:" & " BITSEL_u8_u1_8818_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8818_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8818_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8817_wire_constant, tmp_var);
      BITSEL_u8_u1_8818_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8826_inst flow-through 
    process(BITSEL_u8_u1_8826_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8826_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8825_wire_constant = "& Convert_SLV_To_Hex_String(konst_8825_wire_constant) & " outputs:" & " BITSEL_u8_u1_8826_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8826_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8826_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8825_wire_constant, tmp_var);
      BITSEL_u8_u1_8826_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8834_inst flow-through 
    process(BITSEL_u8_u1_8834_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8834_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8833_wire_constant = "& Convert_SLV_To_Hex_String(konst_8833_wire_constant) & " outputs:" & " BITSEL_u8_u1_8834_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8834_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8834_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8833_wire_constant, tmp_var);
      BITSEL_u8_u1_8834_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8842_inst flow-through 
    process(BITSEL_u8_u1_8842_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8842_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8841_wire_constant = "& Convert_SLV_To_Hex_String(konst_8841_wire_constant) & " outputs:" & " BITSEL_u8_u1_8842_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8842_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8842_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8841_wire_constant, tmp_var);
      BITSEL_u8_u1_8842_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8850_inst flow-through 
    process(BITSEL_u8_u1_8850_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8850_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8849_wire_constant = "& Convert_SLV_To_Hex_String(konst_8849_wire_constant) & " outputs:" & " BITSEL_u8_u1_8850_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8850_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8850_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8849_wire_constant, tmp_var);
      BITSEL_u8_u1_8850_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8858_inst flow-through 
    process(BITSEL_u8_u1_8858_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8858_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8857_wire_constant = "& Convert_SLV_To_Hex_String(konst_8857_wire_constant) & " outputs:" & " BITSEL_u8_u1_8858_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8858_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8858_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8857_wire_constant, tmp_var);
      BITSEL_u8_u1_8858_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8866_inst flow-through 
    process(BITSEL_u8_u1_8866_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8866_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8865_wire_constant = "& Convert_SLV_To_Hex_String(konst_8865_wire_constant) & " outputs:" & " BITSEL_u8_u1_8866_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8866_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8866_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8865_wire_constant, tmp_var);
      BITSEL_u8_u1_8866_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8874_inst flow-through 
    process(BITSEL_u8_u1_8874_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8874_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8873_wire_constant = "& Convert_SLV_To_Hex_String(konst_8873_wire_constant) & " outputs:" & " BITSEL_u8_u1_8874_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8874_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8874_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8873_wire_constant, tmp_var);
      BITSEL_u8_u1_8874_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8882_inst flow-through 
    process(BITSEL_u8_u1_8882_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8882_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8881_wire_constant = "& Convert_SLV_To_Hex_String(konst_8881_wire_constant) & " outputs:" & " BITSEL_u8_u1_8882_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8882_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8882_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8881_wire_constant, tmp_var);
      BITSEL_u8_u1_8882_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8890_inst flow-through 
    process(BITSEL_u8_u1_8890_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8890_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8889_wire_constant = "& Convert_SLV_To_Hex_String(konst_8889_wire_constant) & " outputs:" & " BITSEL_u8_u1_8890_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8890_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8890_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8889_wire_constant, tmp_var);
      BITSEL_u8_u1_8890_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8898_inst flow-through 
    process(BITSEL_u8_u1_8898_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8898_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8897_wire_constant = "& Convert_SLV_To_Hex_String(konst_8897_wire_constant) & " outputs:" & " BITSEL_u8_u1_8898_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8898_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8898_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8897_wire_constant, tmp_var);
      BITSEL_u8_u1_8898_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8906_inst flow-through 
    process(BITSEL_u8_u1_8906_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8906_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8905_wire_constant = "& Convert_SLV_To_Hex_String(konst_8905_wire_constant) & " outputs:" & " BITSEL_u8_u1_8906_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8906_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8906_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8905_wire_constant, tmp_var);
      BITSEL_u8_u1_8906_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8914_inst flow-through 
    process(BITSEL_u8_u1_8914_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8914_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8913_wire_constant = "& Convert_SLV_To_Hex_String(konst_8913_wire_constant) & " outputs:" & " BITSEL_u8_u1_8914_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8914_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8914_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8913_wire_constant, tmp_var);
      BITSEL_u8_u1_8914_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8922_inst flow-through 
    process(BITSEL_u8_u1_8922_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8922_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8921_wire_constant = "& Convert_SLV_To_Hex_String(konst_8921_wire_constant) & " outputs:" & " BITSEL_u8_u1_8922_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8922_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8922_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8921_wire_constant, tmp_var);
      BITSEL_u8_u1_8922_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8930_inst flow-through 
    process(BITSEL_u8_u1_8930_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8930_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8929_wire_constant = "& Convert_SLV_To_Hex_String(konst_8929_wire_constant) & " outputs:" & " BITSEL_u8_u1_8930_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8930_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8930_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8929_wire_constant, tmp_var);
      BITSEL_u8_u1_8930_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8938_inst flow-through 
    process(BITSEL_u8_u1_8938_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8938_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8937_wire_constant = "& Convert_SLV_To_Hex_String(konst_8937_wire_constant) & " outputs:" & " BITSEL_u8_u1_8938_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8938_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8938_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8937_wire_constant, tmp_var);
      BITSEL_u8_u1_8938_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8946_inst flow-through 
    process(BITSEL_u8_u1_8946_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8946_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8945_wire_constant = "& Convert_SLV_To_Hex_String(konst_8945_wire_constant) & " outputs:" & " BITSEL_u8_u1_8946_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8946_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8946_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8945_wire_constant, tmp_var);
      BITSEL_u8_u1_8946_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8954_inst flow-through 
    process(BITSEL_u8_u1_8954_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8954_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8953_wire_constant = "& Convert_SLV_To_Hex_String(konst_8953_wire_constant) & " outputs:" & " BITSEL_u8_u1_8954_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8954_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8954_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8953_wire_constant, tmp_var);
      BITSEL_u8_u1_8954_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8962_inst flow-through 
    process(BITSEL_u8_u1_8962_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8962_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8961_wire_constant = "& Convert_SLV_To_Hex_String(konst_8961_wire_constant) & " outputs:" & " BITSEL_u8_u1_8962_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8962_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8962_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8961_wire_constant, tmp_var);
      BITSEL_u8_u1_8962_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8970_inst flow-through 
    process(BITSEL_u8_u1_8970_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8970_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8969_wire_constant = "& Convert_SLV_To_Hex_String(konst_8969_wire_constant) & " outputs:" & " BITSEL_u8_u1_8970_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8970_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8970_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8969_wire_constant, tmp_var);
      BITSEL_u8_u1_8970_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8978_inst flow-through 
    process(BITSEL_u8_u1_8978_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8978_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8977_wire_constant = "& Convert_SLV_To_Hex_String(konst_8977_wire_constant) & " outputs:" & " BITSEL_u8_u1_8978_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8978_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8978_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8977_wire_constant, tmp_var);
      BITSEL_u8_u1_8978_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8986_inst flow-through 
    process(BITSEL_u8_u1_8986_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8986_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8985_wire_constant = "& Convert_SLV_To_Hex_String(konst_8985_wire_constant) & " outputs:" & " BITSEL_u8_u1_8986_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8986_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8986_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8985_wire_constant, tmp_var);
      BITSEL_u8_u1_8986_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_8994_inst flow-through 
    process(BITSEL_u8_u1_8994_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_8994_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_8993_wire_constant = "& Convert_SLV_To_Hex_String(konst_8993_wire_constant) & " outputs:" & " BITSEL_u8_u1_8994_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_8994_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_8994_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8993_wire_constant, tmp_var);
      BITSEL_u8_u1_8994_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_9002_inst flow-through 
    process(BITSEL_u8_u1_9002_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_9002_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_9001_wire_constant = "& Convert_SLV_To_Hex_String(konst_9001_wire_constant) & " outputs:" & " BITSEL_u8_u1_9002_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_9002_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_9002_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_9001_wire_constant, tmp_var);
      BITSEL_u8_u1_9002_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_9010_inst flow-through 
    process(BITSEL_u8_u1_9010_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_9010_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_9009_wire_constant = "& Convert_SLV_To_Hex_String(konst_9009_wire_constant) & " outputs:" & " BITSEL_u8_u1_9010_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_9010_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_9010_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_9009_wire_constant, tmp_var);
      BITSEL_u8_u1_9010_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_9018_inst flow-through 
    process(BITSEL_u8_u1_9018_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_9018_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_9017_wire_constant = "& Convert_SLV_To_Hex_String(konst_9017_wire_constant) & " outputs:" & " BITSEL_u8_u1_9018_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_9018_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_9018_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_9017_wire_constant, tmp_var);
      BITSEL_u8_u1_9018_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_9026_inst flow-through 
    process(BITSEL_u8_u1_9026_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_9026_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_9025_wire_constant = "& Convert_SLV_To_Hex_String(konst_9025_wire_constant) & " outputs:" & " BITSEL_u8_u1_9026_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_9026_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_9026_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_9025_wire_constant, tmp_var);
      BITSEL_u8_u1_9026_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_9034_inst flow-through 
    process(BITSEL_u8_u1_9034_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_9034_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_9033_wire_constant = "& Convert_SLV_To_Hex_String(konst_9033_wire_constant) & " outputs:" & " BITSEL_u8_u1_9034_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_9034_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_9034_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_9033_wire_constant, tmp_var);
      BITSEL_u8_u1_9034_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_9042_inst flow-through 
    process(BITSEL_u8_u1_9042_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_9042_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_9041_wire_constant = "& Convert_SLV_To_Hex_String(konst_9041_wire_constant) & " outputs:" & " BITSEL_u8_u1_9042_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_9042_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_9042_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_9041_wire_constant, tmp_var);
      BITSEL_u8_u1_9042_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_9050_inst flow-through 
    process(BITSEL_u8_u1_9050_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_9050_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_9049_wire_constant = "& Convert_SLV_To_Hex_String(konst_9049_wire_constant) & " outputs:" & " BITSEL_u8_u1_9050_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_9050_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_9050_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_9049_wire_constant, tmp_var);
      BITSEL_u8_u1_9050_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_9058_inst flow-through 
    process(BITSEL_u8_u1_9058_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_9058_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_9057_wire_constant = "& Convert_SLV_To_Hex_String(konst_9057_wire_constant) & " outputs:" & " BITSEL_u8_u1_9058_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_9058_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_9058_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_9057_wire_constant, tmp_var);
      BITSEL_u8_u1_9058_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_9066_inst flow-through 
    process(BITSEL_u8_u1_9066_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_9066_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_9065_wire_constant = "& Convert_SLV_To_Hex_String(konst_9065_wire_constant) & " outputs:" & " BITSEL_u8_u1_9066_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_9066_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_9066_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_9065_wire_constant, tmp_var);
      BITSEL_u8_u1_9066_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_9074_inst flow-through 
    process(BITSEL_u8_u1_9074_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_9074_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_9073_wire_constant = "& Convert_SLV_To_Hex_String(konst_9073_wire_constant) & " outputs:" & " BITSEL_u8_u1_9074_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_9074_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_9074_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_9073_wire_constant, tmp_var);
      BITSEL_u8_u1_9074_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_9082_inst flow-through 
    process(BITSEL_u8_u1_9082_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_9082_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_9081_wire_constant = "& Convert_SLV_To_Hex_String(konst_9081_wire_constant) & " outputs:" & " BITSEL_u8_u1_9082_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_9082_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_9082_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_9081_wire_constant, tmp_var);
      BITSEL_u8_u1_9082_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_9090_inst flow-through 
    process(BITSEL_u8_u1_9090_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_9090_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_9089_wire_constant = "& Convert_SLV_To_Hex_String(konst_9089_wire_constant) & " outputs:" & " BITSEL_u8_u1_9090_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_9090_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_9090_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_9089_wire_constant, tmp_var);
      BITSEL_u8_u1_9090_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_9098_inst flow-through 
    process(BITSEL_u8_u1_9098_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_9098_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_9097_wire_constant = "& Convert_SLV_To_Hex_String(konst_9097_wire_constant) & " outputs:" & " BITSEL_u8_u1_9098_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_9098_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_9098_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_9097_wire_constant, tmp_var);
      BITSEL_u8_u1_9098_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_9106_inst flow-through 
    process(BITSEL_u8_u1_9106_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_9106_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_9105_wire_constant = "& Convert_SLV_To_Hex_String(konst_9105_wire_constant) & " outputs:" & " BITSEL_u8_u1_9106_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_9106_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_9106_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_9105_wire_constant, tmp_var);
      BITSEL_u8_u1_9106_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_9114_inst flow-through 
    process(BITSEL_u8_u1_9114_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_9114_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_9113_wire_constant = "& Convert_SLV_To_Hex_String(konst_9113_wire_constant) & " outputs:" & " BITSEL_u8_u1_9114_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_9114_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_9114_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_9113_wire_constant, tmp_var);
      BITSEL_u8_u1_9114_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_9122_inst flow-through 
    process(BITSEL_u8_u1_9122_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_9122_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_9121_wire_constant = "& Convert_SLV_To_Hex_String(konst_9121_wire_constant) & " outputs:" & " BITSEL_u8_u1_9122_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_9122_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_9122_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_9121_wire_constant, tmp_var);
      BITSEL_u8_u1_9122_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_9130_inst flow-through 
    process(BITSEL_u8_u1_9130_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_9130_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_9129_wire_constant = "& Convert_SLV_To_Hex_String(konst_9129_wire_constant) & " outputs:" & " BITSEL_u8_u1_9130_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_9130_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_9130_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_9129_wire_constant, tmp_var);
      BITSEL_u8_u1_9130_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_9138_inst flow-through 
    process(BITSEL_u8_u1_9138_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_9138_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_9137_wire_constant = "& Convert_SLV_To_Hex_String(konst_9137_wire_constant) & " outputs:" & " BITSEL_u8_u1_9138_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_9138_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_9138_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_9137_wire_constant, tmp_var);
      BITSEL_u8_u1_9138_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_9146_inst flow-through 
    process(BITSEL_u8_u1_9146_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_9146_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_9145_wire_constant = "& Convert_SLV_To_Hex_String(konst_9145_wire_constant) & " outputs:" & " BITSEL_u8_u1_9146_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_9146_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_9146_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_9145_wire_constant, tmp_var);
      BITSEL_u8_u1_9146_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_9154_inst flow-through 
    process(BITSEL_u8_u1_9154_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_9154_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_9153_wire_constant = "& Convert_SLV_To_Hex_String(konst_9153_wire_constant) & " outputs:" & " BITSEL_u8_u1_9154_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_9154_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_9154_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_9153_wire_constant, tmp_var);
      BITSEL_u8_u1_9154_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_9162_inst flow-through 
    process(BITSEL_u8_u1_9162_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_9162_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_9161_wire_constant = "& Convert_SLV_To_Hex_String(konst_9161_wire_constant) & " outputs:" & " BITSEL_u8_u1_9162_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_9162_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_9162_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_9161_wire_constant, tmp_var);
      BITSEL_u8_u1_9162_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_9170_inst flow-through 
    process(BITSEL_u8_u1_9170_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_9170_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_9169_wire_constant = "& Convert_SLV_To_Hex_String(konst_9169_wire_constant) & " outputs:" & " BITSEL_u8_u1_9170_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_9170_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_9170_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_9169_wire_constant, tmp_var);
      BITSEL_u8_u1_9170_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_9178_inst flow-through 
    process(BITSEL_u8_u1_9178_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_9178_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_9177_wire_constant = "& Convert_SLV_To_Hex_String(konst_9177_wire_constant) & " outputs:" & " BITSEL_u8_u1_9178_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_9178_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_9178_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_9177_wire_constant, tmp_var);
      BITSEL_u8_u1_9178_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_9186_inst flow-through 
    process(BITSEL_u8_u1_9186_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_9186_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_9185_wire_constant = "& Convert_SLV_To_Hex_String(konst_9185_wire_constant) & " outputs:" & " BITSEL_u8_u1_9186_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_9186_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_9186_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_9185_wire_constant, tmp_var);
      BITSEL_u8_u1_9186_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_9194_inst flow-through 
    process(BITSEL_u8_u1_9194_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_9194_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_9193_wire_constant = "& Convert_SLV_To_Hex_String(konst_9193_wire_constant) & " outputs:" & " BITSEL_u8_u1_9194_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_9194_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_9194_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_9193_wire_constant, tmp_var);
      BITSEL_u8_u1_9194_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator BITSEL_u8_u1_9202_inst flow-through 
    process(BITSEL_u8_u1_9202_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:Inv_Sbox_4:DP:BITSEL_u8_u1_9202_inst:flowthrough inputs: " & " s_in_buffer = "& Convert_SLV_To_Hex_String(s_in_buffer) & " konst_9201_wire_constant = "& Convert_SLV_To_Hex_String(konst_9201_wire_constant) & " outputs:" & " BITSEL_u8_u1_9202_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_9202_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_9202_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_9201_wire_constant, tmp_var);
      BITSEL_u8_u1_9202_wire <= tmp_var; -- 
    end process;
    -- 
  end Block; -- data_path
  -- 
end Inv_Sbox_4_Volatile_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library GhdlLink;
use GhdlLink.LogUtilities.all;
library work;
use work.ahir_system_global_package.all;
entity MUL2_Volatile is -- 
  port ( -- 
    clk, reset: in std_logic; 
    mul_in : in  std_logic_vector(7 downto 0);
    mul_out : out  std_logic_vector(7 downto 0)-- 
  );
  -- 
end entity MUL2_Volatile;
architecture MUL2_Volatile_arch of MUL2_Volatile is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector(8-1 downto 0);
  signal default_zero_sig: std_logic;
  -- input port buffer signals
  signal mul_in_buffer :  std_logic_vector(7 downto 0);
  -- output port buffer signals
  signal mul_out_buffer :  std_logic_vector(7 downto 0);
  -- volatile/operator module components. 
  signal global_clock_cycle_count: integer := 0;
  -- 
begin --  
  ---------------------------------------------------------- 
  process(clk)  
  begin -- 
    if(clk'event and clk = '1') then -- 
      if(reset = '1') then -- 
        global_clock_cycle_count <= 0; --
      else -- 
        global_clock_cycle_count <= global_clock_cycle_count + 1; -- 
      end if; --
    end if; --
  end process;
  ---------------------------------------------------------- 
  -- input handling ------------------------------------------------
  mul_in_buffer <= mul_in;
  -- output handling  -------------------------------------------------------
  mul_out <= mul_out_buffer;
  -- the control path --------------------------------------------------
  default_zero_sig <= '0';
  -- volatile module, no control path
  -- the data path
  data_path: Block -- 
    signal BITSEL_u8_u1_9222_wire : std_logic_vector(0 downto 0);
    signal R_mod_const_9224_wire_constant : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_9225_wire : std_logic_vector(7 downto 0);
    signal inx2_9218 : std_logic_vector(7 downto 0);
    signal konst_9216_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9221_wire_constant : std_logic_vector(7 downto 0);
    signal xxMUL2xxmod_const : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    R_mod_const_9224_wire_constant <= "00011011";
    konst_9216_wire_constant <= "00000001";
    konst_9221_wire_constant <= "00000111";
    xxMUL2xxmod_const <= "00011011";
    -- logger for split-operator MUX_9227_inst flow-through 
    process(mul_out_buffer) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:MUL2:DP:MUX_9227_inst:flowthrough inputs: " & " BITSEL_u8_u1_9222_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_9222_wire) & " XOR_u8_u8_9225_wire = "& Convert_SLV_To_Hex_String(XOR_u8_u8_9225_wire) & " inx2_9218 = "& Convert_SLV_To_Hex_String(inx2_9218) & " outputs:" & " mul_out_buffer= "  & Convert_SLV_To_Hex_String(mul_out_buffer));
      --
    end process; 
    -- flow-through select operator MUX_9227_inst
    mul_out_buffer <= XOR_u8_u8_9225_wire when (BITSEL_u8_u1_9222_wire(0) /=  '0') else inx2_9218;
    -- logger for split-operator BITSEL_u8_u1_9222_inst flow-through 
    process(BITSEL_u8_u1_9222_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:MUL2:DP:BITSEL_u8_u1_9222_inst:flowthrough inputs: " & " mul_in_buffer = "& Convert_SLV_To_Hex_String(mul_in_buffer) & " konst_9221_wire_constant = "& Convert_SLV_To_Hex_String(konst_9221_wire_constant) & " outputs:" & " BITSEL_u8_u1_9222_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_9222_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_9222_inst
    process(mul_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(mul_in_buffer, konst_9221_wire_constant, tmp_var);
      BITSEL_u8_u1_9222_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator SHL_u8_u8_9217_inst flow-through 
    process(inx2_9218) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:MUL2:DP:SHL_u8_u8_9217_inst:flowthrough inputs: " & " mul_in_buffer = "& Convert_SLV_To_Hex_String(mul_in_buffer) & " konst_9216_wire_constant = "& Convert_SLV_To_Hex_String(konst_9216_wire_constant) & " outputs:" & " inx2_9218= "  & Convert_SLV_To_Hex_String(inx2_9218));
      --
    end process; 
    -- binary operator SHL_u8_u8_9217_inst
    process(mul_in_buffer) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntSHL_proc(mul_in_buffer, konst_9216_wire_constant, tmp_var);
      inx2_9218 <= tmp_var; -- 
    end process;
    -- logger for split-operator XOR_u8_u8_9225_inst flow-through 
    process(XOR_u8_u8_9225_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:MUL2:DP:XOR_u8_u8_9225_inst:flowthrough inputs: " & " inx2_9218 = "& Convert_SLV_To_Hex_String(inx2_9218) & " R_mod_const_9224_wire_constant = "& Convert_SLV_To_Hex_String(R_mod_const_9224_wire_constant) & " outputs:" & " XOR_u8_u8_9225_wire= "  & Convert_SLV_To_Hex_String(XOR_u8_u8_9225_wire));
      --
    end process; 
    -- binary operator XOR_u8_u8_9225_inst
    process(inx2_9218) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(inx2_9218, R_mod_const_9224_wire_constant, tmp_var);
      XOR_u8_u8_9225_wire <= tmp_var; -- 
    end process;
    -- 
  end Block; -- data_path
  -- 
end MUL2_Volatile_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library GhdlLink;
use GhdlLink.LogUtilities.all;
library work;
use work.ahir_system_global_package.all;
entity c_block_daemon_in is -- 
  generic (tag_length : integer); 
  port ( -- 
    in_data_pipe_read_req : out  std_logic_vector(0 downto 0);
    in_data_pipe_read_ack : in   std_logic_vector(0 downto 0);
    in_data_pipe_read_data : in   std_logic_vector(63 downto 0);
    in_buf_pipe_write_req : out  std_logic_vector(0 downto 0);
    in_buf_pipe_write_ack : in   std_logic_vector(0 downto 0);
    in_buf_pipe_write_data : out  std_logic_vector(127 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity c_block_daemon_in;
architecture c_block_daemon_in_arch of c_block_daemon_in is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal c_block_daemon_in_CP_15_start: Boolean;
  signal c_block_daemon_in_CP_15_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal RPIPE_in_data_9232_inst_req_0 : boolean;
  signal RPIPE_in_data_9232_inst_ack_0 : boolean;
  signal RPIPE_in_data_9232_inst_req_1 : boolean;
  signal RPIPE_in_data_9232_inst_ack_1 : boolean;
  signal RPIPE_in_data_9235_inst_req_0 : boolean;
  signal RPIPE_in_data_9235_inst_ack_0 : boolean;
  signal RPIPE_in_data_9235_inst_req_1 : boolean;
  signal RPIPE_in_data_9235_inst_ack_1 : boolean;
  signal CONCAT_u64_u128_9240_inst_req_0 : boolean;
  signal CONCAT_u64_u128_9240_inst_ack_0 : boolean;
  signal CONCAT_u64_u128_9240_inst_req_1 : boolean;
  signal CONCAT_u64_u128_9240_inst_ack_1 : boolean;
  signal WPIPE_in_buf_9237_inst_req_0 : boolean;
  signal WPIPE_in_buf_9237_inst_ack_0 : boolean;
  signal WPIPE_in_buf_9237_inst_req_1 : boolean;
  signal WPIPE_in_buf_9237_inst_ack_1 : boolean;
  signal global_clock_cycle_count: integer := 0;
  -- 
begin --  
  ---------------------------------------------------------- 
  process(clk)  
  begin -- 
    if(clk'event and clk = '1') then -- 
      if(reset = '1') then -- 
        global_clock_cycle_count <= 0; --
      else -- 
        global_clock_cycle_count <= global_clock_cycle_count + 1; -- 
      end if; --
    end if; --
  end process;
  ---------------------------------------------------------- 
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "c_block_daemon_in_input_buffer", -- 
      buffer_size => 1,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  c_block_daemon_in_CP_15_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "c_block_daemon_in_out_buffer", -- 
      buffer_size => 1,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= c_block_daemon_in_CP_15_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= c_block_daemon_in_CP_15_start & tag_ilock_write_ack_symbol;
    gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= c_block_daemon_in_CP_15_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  --- logging ------------------------------------------------------
  LogCPEvent(clk,reset,global_clock_cycle_count,c_block_daemon_in_CP_15_start,"c_block_daemon_in cp_entry_symbol ");
  LogCPEvent(clk,reset,global_clock_cycle_count,c_block_daemon_in_CP_15_symbol, "c_block_daemon_in cp_exit_symbol ");
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  c_block_daemon_in_CP_15: Block -- control-path 
    signal c_block_daemon_in_CP_15_elements: BooleanArray(8 downto 0);
    -- 
  begin -- 
    c_block_daemon_in_CP_15_elements(0) <= c_block_daemon_in_CP_15_start;
    c_block_daemon_in_CP_15_symbol <= c_block_daemon_in_CP_15_elements(8);
    -- CP-element group 0:  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (5) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_9233/$entry
      -- CP-element group 0: 	 assign_stmt_9233/RPIPE_in_data_9232_sample_start_
      -- CP-element group 0: 	 assign_stmt_9233/RPIPE_in_data_9232_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9233/RPIPE_in_data_9232_Sample/rr
      -- 
    -- logger for CP element group c_block_daemon_in_CP_15_elements(0)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and c_block_daemon_in_CP_15_elements(0)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:c_block_daemon_in:CP:c_block_daemon_in_CP_15_elements(0) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:c_block_daemon_in:CP:RPIPE_in_data_9232_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_28_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => c_block_daemon_in_CP_15_elements(0), ack => RPIPE_in_data_9232_inst_req_0); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 assign_stmt_9233/RPIPE_in_data_9232_sample_completed_
      -- CP-element group 1: 	 assign_stmt_9233/RPIPE_in_data_9232_update_start_
      -- CP-element group 1: 	 assign_stmt_9233/RPIPE_in_data_9232_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_9233/RPIPE_in_data_9232_Sample/ra
      -- CP-element group 1: 	 assign_stmt_9233/RPIPE_in_data_9232_Update/$entry
      -- CP-element group 1: 	 assign_stmt_9233/RPIPE_in_data_9232_Update/cr
      -- 
    -- logger for CP element group c_block_daemon_in_CP_15_elements(1)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and c_block_daemon_in_CP_15_elements(1)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:c_block_daemon_in:CP:c_block_daemon_in_CP_15_elements(1) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:c_block_daemon_in:CP:RPIPE_in_data_9232_inst_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:c_block_daemon_in:CP:RPIPE_in_data_9232_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ra_29_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_in_data_9232_inst_ack_0, ack => c_block_daemon_in_CP_15_elements(1)); -- 
    cr_33_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => c_block_daemon_in_CP_15_elements(1), ack => RPIPE_in_data_9232_inst_req_1); -- 
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (8) 
      -- CP-element group 2: 	 assign_stmt_9233/$exit
      -- CP-element group 2: 	 assign_stmt_9233/RPIPE_in_data_9232_update_completed_
      -- CP-element group 2: 	 assign_stmt_9233/RPIPE_in_data_9232_Update/$exit
      -- CP-element group 2: 	 assign_stmt_9233/RPIPE_in_data_9232_Update/ca
      -- CP-element group 2: 	 assign_stmt_9236/$entry
      -- CP-element group 2: 	 assign_stmt_9236/RPIPE_in_data_9235_sample_start_
      -- CP-element group 2: 	 assign_stmt_9236/RPIPE_in_data_9235_Sample/$entry
      -- CP-element group 2: 	 assign_stmt_9236/RPIPE_in_data_9235_Sample/rr
      -- 
    -- logger for CP element group c_block_daemon_in_CP_15_elements(2)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and c_block_daemon_in_CP_15_elements(2)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:c_block_daemon_in:CP:c_block_daemon_in_CP_15_elements(2) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:c_block_daemon_in:CP:RPIPE_in_data_9232_inst_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:c_block_daemon_in:CP:RPIPE_in_data_9235_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ca_34_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_in_data_9232_inst_ack_1, ack => c_block_daemon_in_CP_15_elements(2)); -- 
    rr_45_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => c_block_daemon_in_CP_15_elements(2), ack => RPIPE_in_data_9235_inst_req_0); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 assign_stmt_9236/RPIPE_in_data_9235_sample_completed_
      -- CP-element group 3: 	 assign_stmt_9236/RPIPE_in_data_9235_update_start_
      -- CP-element group 3: 	 assign_stmt_9236/RPIPE_in_data_9235_Sample/$exit
      -- CP-element group 3: 	 assign_stmt_9236/RPIPE_in_data_9235_Sample/ra
      -- CP-element group 3: 	 assign_stmt_9236/RPIPE_in_data_9235_Update/$entry
      -- CP-element group 3: 	 assign_stmt_9236/RPIPE_in_data_9235_Update/cr
      -- 
    -- logger for CP element group c_block_daemon_in_CP_15_elements(3)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and c_block_daemon_in_CP_15_elements(3)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:c_block_daemon_in:CP:c_block_daemon_in_CP_15_elements(3) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:c_block_daemon_in:CP:RPIPE_in_data_9235_inst_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:c_block_daemon_in:CP:RPIPE_in_data_9235_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ra_46_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_in_data_9235_inst_ack_0, ack => c_block_daemon_in_CP_15_elements(3)); -- 
    cr_50_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => c_block_daemon_in_CP_15_elements(3), ack => RPIPE_in_data_9235_inst_req_1); -- 
    -- CP-element group 4:  join  fork  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	6 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (19) 
      -- CP-element group 4: 	 assign_stmt_9236/$exit
      -- CP-element group 4: 	 assign_stmt_9236/RPIPE_in_data_9235_update_completed_
      -- CP-element group 4: 	 assign_stmt_9236/RPIPE_in_data_9235_Update/$exit
      -- CP-element group 4: 	 assign_stmt_9236/RPIPE_in_data_9235_Update/ca
      -- CP-element group 4: 	 assign_stmt_9241/$entry
      -- CP-element group 4: 	 assign_stmt_9241/CONCAT_u64_u128_9240_sample_start_
      -- CP-element group 4: 	 assign_stmt_9241/CONCAT_u64_u128_9240_update_start_
      -- CP-element group 4: 	 assign_stmt_9241/R_Ina_9238_sample_start_
      -- CP-element group 4: 	 assign_stmt_9241/R_Ina_9238_sample_completed_
      -- CP-element group 4: 	 assign_stmt_9241/R_Ina_9238_update_start_
      -- CP-element group 4: 	 assign_stmt_9241/R_Ina_9238_update_completed_
      -- CP-element group 4: 	 assign_stmt_9241/R_Inb_9239_sample_start_
      -- CP-element group 4: 	 assign_stmt_9241/R_Inb_9239_sample_completed_
      -- CP-element group 4: 	 assign_stmt_9241/R_Inb_9239_update_start_
      -- CP-element group 4: 	 assign_stmt_9241/R_Inb_9239_update_completed_
      -- CP-element group 4: 	 assign_stmt_9241/CONCAT_u64_u128_9240_Sample/$entry
      -- CP-element group 4: 	 assign_stmt_9241/CONCAT_u64_u128_9240_Sample/rr
      -- CP-element group 4: 	 assign_stmt_9241/CONCAT_u64_u128_9240_Update/$entry
      -- CP-element group 4: 	 assign_stmt_9241/CONCAT_u64_u128_9240_Update/cr
      -- 
    -- logger for CP element group c_block_daemon_in_CP_15_elements(4)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and c_block_daemon_in_CP_15_elements(4)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:c_block_daemon_in:CP:c_block_daemon_in_CP_15_elements(4) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:c_block_daemon_in:CP:RPIPE_in_data_9235_inst_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:c_block_daemon_in:CP:CONCAT_u64_u128_9240_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:c_block_daemon_in:CP:CONCAT_u64_u128_9240_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ca_51_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_in_data_9235_inst_ack_1, ack => c_block_daemon_in_CP_15_elements(4)); -- 
    cr_75_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => c_block_daemon_in_CP_15_elements(4), ack => CONCAT_u64_u128_9240_inst_req_1); -- 
    rr_70_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => c_block_daemon_in_CP_15_elements(4), ack => CONCAT_u64_u128_9240_inst_req_0); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 assign_stmt_9241/CONCAT_u64_u128_9240_sample_completed_
      -- CP-element group 5: 	 assign_stmt_9241/CONCAT_u64_u128_9240_Sample/$exit
      -- CP-element group 5: 	 assign_stmt_9241/CONCAT_u64_u128_9240_Sample/ra
      -- 
    -- logger for CP element group c_block_daemon_in_CP_15_elements(5)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and c_block_daemon_in_CP_15_elements(5)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:c_block_daemon_in:CP:c_block_daemon_in_CP_15_elements(5) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:c_block_daemon_in:CP:CONCAT_u64_u128_9240_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_71_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u64_u128_9240_inst_ack_0, ack => c_block_daemon_in_CP_15_elements(5)); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	4 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (6) 
      -- CP-element group 6: 	 assign_stmt_9241/CONCAT_u64_u128_9240_update_completed_
      -- CP-element group 6: 	 assign_stmt_9241/CONCAT_u64_u128_9240_Update/$exit
      -- CP-element group 6: 	 assign_stmt_9241/CONCAT_u64_u128_9240_Update/ca
      -- CP-element group 6: 	 assign_stmt_9241/WPIPE_in_buf_9237_sample_start_
      -- CP-element group 6: 	 assign_stmt_9241/WPIPE_in_buf_9237_Sample/$entry
      -- CP-element group 6: 	 assign_stmt_9241/WPIPE_in_buf_9237_Sample/req
      -- 
    -- logger for CP element group c_block_daemon_in_CP_15_elements(6)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and c_block_daemon_in_CP_15_elements(6)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:c_block_daemon_in:CP:c_block_daemon_in_CP_15_elements(6) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:c_block_daemon_in:CP:CONCAT_u64_u128_9240_inst_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:c_block_daemon_in:CP:WPIPE_in_buf_9237_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ca_76_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u64_u128_9240_inst_ack_1, ack => c_block_daemon_in_CP_15_elements(6)); -- 
    req_84_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => c_block_daemon_in_CP_15_elements(6), ack => WPIPE_in_buf_9237_inst_req_0); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 assign_stmt_9241/WPIPE_in_buf_9237_sample_completed_
      -- CP-element group 7: 	 assign_stmt_9241/WPIPE_in_buf_9237_update_start_
      -- CP-element group 7: 	 assign_stmt_9241/WPIPE_in_buf_9237_Sample/$exit
      -- CP-element group 7: 	 assign_stmt_9241/WPIPE_in_buf_9237_Sample/ack
      -- CP-element group 7: 	 assign_stmt_9241/WPIPE_in_buf_9237_Update/$entry
      -- CP-element group 7: 	 assign_stmt_9241/WPIPE_in_buf_9237_Update/req
      -- 
    -- logger for CP element group c_block_daemon_in_CP_15_elements(7)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and c_block_daemon_in_CP_15_elements(7)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:c_block_daemon_in:CP:c_block_daemon_in_CP_15_elements(7) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:c_block_daemon_in:CP:WPIPE_in_buf_9237_inst_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:c_block_daemon_in:CP:WPIPE_in_buf_9237_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_85_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_in_buf_9237_inst_ack_0, ack => c_block_daemon_in_CP_15_elements(7)); -- 
    req_89_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => c_block_daemon_in_CP_15_elements(7), ack => WPIPE_in_buf_9237_inst_req_1); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8:  members (5) 
      -- CP-element group 8: 	 $exit
      -- CP-element group 8: 	 assign_stmt_9241/$exit
      -- CP-element group 8: 	 assign_stmt_9241/WPIPE_in_buf_9237_update_completed_
      -- CP-element group 8: 	 assign_stmt_9241/WPIPE_in_buf_9237_Update/$exit
      -- CP-element group 8: 	 assign_stmt_9241/WPIPE_in_buf_9237_Update/ack
      -- 
    -- logger for CP element group c_block_daemon_in_CP_15_elements(8)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and c_block_daemon_in_CP_15_elements(8)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:c_block_daemon_in:CP:c_block_daemon_in_CP_15_elements(8) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:c_block_daemon_in:CP:WPIPE_in_buf_9237_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_90_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_in_buf_9237_inst_ack_1, ack => c_block_daemon_in_CP_15_elements(8)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal CONCAT_u64_u128_9240_wire : std_logic_vector(127 downto 0);
    signal Ina_9233 : std_logic_vector(63 downto 0);
    signal Inb_9236 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    -- logger for split-operator CONCAT_u64_u128_9240_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if CONCAT_u64_u128_9240_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:c_block_daemon_in:DP:CONCAT_u64_u128_9240_inst:started:   inputs: " & " Ina_9233 = "& Convert_SLV_To_Hex_String(Ina_9233) & " Inb_9236 = "& Convert_SLV_To_Hex_String(Inb_9236));
          --
        end if; 
        if CONCAT_u64_u128_9240_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:c_block_daemon_in:DP:CONCAT_u64_u128_9240_inst:finished:  outputs: " & " CONCAT_u64_u128_9240_wire= "  & Convert_SLV_To_Hex_String(CONCAT_u64_u128_9240_wire));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (0) : CONCAT_u64_u128_9240_inst 
    ApConcat_group_0: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= Ina_9233 & Inb_9236;
      CONCAT_u64_u128_9240_wire <= data_out(127 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= CONCAT_u64_u128_9240_inst_req_0;
      CONCAT_u64_u128_9240_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= CONCAT_u64_u128_9240_inst_req_1;
      CONCAT_u64_u128_9240_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApConcat",
          name => "ApConcat_group_0",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 64, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 128,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- logger for split-operator RPIPE_in_data_9232_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if RPIPE_in_data_9232_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:c_block_daemon_in:DP:RPIPE_in_data_9232_inst:started:   PipeRead from in_data inputs: " & " no-guard, no-inputs ");
          --
        end if; 
        if RPIPE_in_data_9232_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:c_block_daemon_in:DP:RPIPE_in_data_9232_inst:finished:  outputs: " & " Ina_9233= "  & Convert_SLV_To_Hex_String(Ina_9233));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator RPIPE_in_data_9235_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if RPIPE_in_data_9235_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:c_block_daemon_in:DP:RPIPE_in_data_9235_inst:started:   PipeRead from in_data inputs: " & " no-guard, no-inputs ");
          --
        end if; 
        if RPIPE_in_data_9235_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:c_block_daemon_in:DP:RPIPE_in_data_9235_inst:finished:  outputs: " & " Inb_9236= "  & Convert_SLV_To_Hex_String(Inb_9236));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared inport operator group (0) : RPIPE_in_data_9232_inst RPIPE_in_data_9235_inst 
    InportGroup0: Block -- 
      signal data_out: std_logic_vector(127 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 1 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= RPIPE_in_data_9232_inst_req_0;
      reqL_unguarded(0) <= RPIPE_in_data_9235_inst_req_0;
      RPIPE_in_data_9232_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_in_data_9235_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= RPIPE_in_data_9232_inst_req_1;
      reqR_unguarded(0) <= RPIPE_in_data_9235_inst_req_1;
      RPIPE_in_data_9232_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_in_data_9235_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      gI: SplitGuardInterface generic map(nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Ina_9233 <= data_out(127 downto 64);
      Inb_9236 <= data_out(63 downto 0);
      in_data_read_0: InputPortRevised -- 
        generic map ( name => "in_data_read_0", data_width => 64,  num_reqs => 2,  output_buffering => outBUFs,   no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => in_data_pipe_read_req(0),
          oack => in_data_pipe_read_ack(0),
          odata => in_data_pipe_read_data(63 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- logger for split-operator WPIPE_in_buf_9237_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if WPIPE_in_buf_9237_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:c_block_daemon_in:DP:WPIPE_in_buf_9237_inst:started:   PipeWrite to in_buf inputs: " & " CONCAT_u64_u128_9240_wire = "& Convert_SLV_To_Hex_String(CONCAT_u64_u128_9240_wire));
          --
        end if; 
        if WPIPE_in_buf_9237_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:c_block_daemon_in:DP:WPIPE_in_buf_9237_inst:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared outport operator group (0) : WPIPE_in_buf_9237_inst 
    OutportGroup0: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_in_buf_9237_inst_req_0;
      WPIPE_in_buf_9237_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_in_buf_9237_inst_req_1;
      WPIPE_in_buf_9237_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      data_in <= CONCAT_u64_u128_9240_wire;
      in_buf_write_0: OutputPortRevised -- 
        generic map ( name => "in_buf", data_width => 128, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => in_buf_pipe_write_req(0),
          oack => in_buf_pipe_write_ack(0),
          odata => in_buf_pipe_write_data(127 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end c_block_daemon_in_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library GhdlLink;
use GhdlLink.LogUtilities.all;
library work;
use work.ahir_system_global_package.all;
entity c_block_daemon_out is -- 
  generic (tag_length : integer); 
  port ( -- 
    out_buf_pipe_read_req : out  std_logic_vector(0 downto 0);
    out_buf_pipe_read_ack : in   std_logic_vector(0 downto 0);
    out_buf_pipe_read_data : in   std_logic_vector(127 downto 0);
    out_data_pipe_write_req : out  std_logic_vector(0 downto 0);
    out_data_pipe_write_ack : in   std_logic_vector(0 downto 0);
    out_data_pipe_write_data : out  std_logic_vector(63 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity c_block_daemon_out;
architecture c_block_daemon_out_arch of c_block_daemon_out is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal c_block_daemon_out_CP_91_start: Boolean;
  signal c_block_daemon_out_CP_91_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal RPIPE_out_buf_9245_inst_req_0 : boolean;
  signal RPIPE_out_buf_9245_inst_ack_0 : boolean;
  signal RPIPE_out_buf_9245_inst_req_1 : boolean;
  signal RPIPE_out_buf_9245_inst_ack_1 : boolean;
  signal WPIPE_out_data_9255_inst_req_0 : boolean;
  signal WPIPE_out_data_9255_inst_ack_0 : boolean;
  signal WPIPE_out_data_9255_inst_req_1 : boolean;
  signal WPIPE_out_data_9255_inst_ack_1 : boolean;
  signal WPIPE_out_data_9258_inst_req_0 : boolean;
  signal WPIPE_out_data_9258_inst_ack_0 : boolean;
  signal WPIPE_out_data_9258_inst_req_1 : boolean;
  signal WPIPE_out_data_9258_inst_ack_1 : boolean;
  signal global_clock_cycle_count: integer := 0;
  -- 
begin --  
  ---------------------------------------------------------- 
  process(clk)  
  begin -- 
    if(clk'event and clk = '1') then -- 
      if(reset = '1') then -- 
        global_clock_cycle_count <= 0; --
      else -- 
        global_clock_cycle_count <= global_clock_cycle_count + 1; -- 
      end if; --
    end if; --
  end process;
  ---------------------------------------------------------- 
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "c_block_daemon_out_input_buffer", -- 
      buffer_size => 1,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  c_block_daemon_out_CP_91_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "c_block_daemon_out_out_buffer", -- 
      buffer_size => 1,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= c_block_daemon_out_CP_91_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= c_block_daemon_out_CP_91_start & tag_ilock_write_ack_symbol;
    gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= c_block_daemon_out_CP_91_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  --- logging ------------------------------------------------------
  LogCPEvent(clk,reset,global_clock_cycle_count,c_block_daemon_out_CP_91_start,"c_block_daemon_out cp_entry_symbol ");
  LogCPEvent(clk,reset,global_clock_cycle_count,c_block_daemon_out_CP_91_symbol, "c_block_daemon_out cp_exit_symbol ");
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  c_block_daemon_out_CP_91: Block -- control-path 
    signal c_block_daemon_out_CP_91_elements: BooleanArray(6 downto 0);
    -- 
  begin -- 
    c_block_daemon_out_CP_91_elements(0) <= c_block_daemon_out_CP_91_start;
    c_block_daemon_out_CP_91_symbol <= c_block_daemon_out_CP_91_elements(6);
    -- CP-element group 0:  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (5) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_9246/$entry
      -- CP-element group 0: 	 assign_stmt_9246/RPIPE_out_buf_9245_sample_start_
      -- CP-element group 0: 	 assign_stmt_9246/RPIPE_out_buf_9245_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9246/RPIPE_out_buf_9245_Sample/rr
      -- 
    -- logger for CP element group c_block_daemon_out_CP_91_elements(0)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and c_block_daemon_out_CP_91_elements(0)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:c_block_daemon_out:CP:c_block_daemon_out_CP_91_elements(0) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:c_block_daemon_out:CP:RPIPE_out_buf_9245_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_104_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => c_block_daemon_out_CP_91_elements(0), ack => RPIPE_out_buf_9245_inst_req_0); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 assign_stmt_9246/RPIPE_out_buf_9245_sample_completed_
      -- CP-element group 1: 	 assign_stmt_9246/RPIPE_out_buf_9245_update_start_
      -- CP-element group 1: 	 assign_stmt_9246/RPIPE_out_buf_9245_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_9246/RPIPE_out_buf_9245_Sample/ra
      -- CP-element group 1: 	 assign_stmt_9246/RPIPE_out_buf_9245_Update/$entry
      -- CP-element group 1: 	 assign_stmt_9246/RPIPE_out_buf_9245_Update/cr
      -- 
    -- logger for CP element group c_block_daemon_out_CP_91_elements(1)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and c_block_daemon_out_CP_91_elements(1)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:c_block_daemon_out:CP:c_block_daemon_out_CP_91_elements(1) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:c_block_daemon_out:CP:RPIPE_out_buf_9245_inst_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:c_block_daemon_out:CP:RPIPE_out_buf_9245_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ra_105_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_out_buf_9245_inst_ack_0, ack => c_block_daemon_out_CP_91_elements(1)); -- 
    cr_109_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => c_block_daemon_out_CP_91_elements(1), ack => RPIPE_out_buf_9245_inst_req_1); -- 
    -- CP-element group 2:  join  fork  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (46) 
      -- CP-element group 2: 	 assign_stmt_9246/$exit
      -- CP-element group 2: 	 assign_stmt_9246/RPIPE_out_buf_9245_update_completed_
      -- CP-element group 2: 	 assign_stmt_9246/RPIPE_out_buf_9245_Update/$exit
      -- CP-element group 2: 	 assign_stmt_9246/RPIPE_out_buf_9245_Update/ca
      -- CP-element group 2: 	 assign_stmt_9250_to_assign_stmt_9254/$entry
      -- CP-element group 2: 	 assign_stmt_9250_to_assign_stmt_9254/$exit
      -- CP-element group 2: 	 assign_stmt_9250_to_assign_stmt_9254/slice_9249_sample_start_
      -- CP-element group 2: 	 assign_stmt_9250_to_assign_stmt_9254/slice_9249_sample_completed_
      -- CP-element group 2: 	 assign_stmt_9250_to_assign_stmt_9254/slice_9249_update_start_
      -- CP-element group 2: 	 assign_stmt_9250_to_assign_stmt_9254/slice_9249_update_completed_
      -- CP-element group 2: 	 assign_stmt_9250_to_assign_stmt_9254/R_Z_9248_sample_start_
      -- CP-element group 2: 	 assign_stmt_9250_to_assign_stmt_9254/R_Z_9248_sample_completed_
      -- CP-element group 2: 	 assign_stmt_9250_to_assign_stmt_9254/R_Z_9248_update_start_
      -- CP-element group 2: 	 assign_stmt_9250_to_assign_stmt_9254/R_Z_9248_update_completed_
      -- CP-element group 2: 	 assign_stmt_9250_to_assign_stmt_9254/slice_9249_Sample/$entry
      -- CP-element group 2: 	 assign_stmt_9250_to_assign_stmt_9254/slice_9249_Sample/$exit
      -- CP-element group 2: 	 assign_stmt_9250_to_assign_stmt_9254/slice_9249_Sample/rr
      -- CP-element group 2: 	 assign_stmt_9250_to_assign_stmt_9254/slice_9249_Sample/ra
      -- CP-element group 2: 	 assign_stmt_9250_to_assign_stmt_9254/slice_9249_Update/$entry
      -- CP-element group 2: 	 assign_stmt_9250_to_assign_stmt_9254/slice_9249_Update/$exit
      -- CP-element group 2: 	 assign_stmt_9250_to_assign_stmt_9254/slice_9249_Update/cr
      -- CP-element group 2: 	 assign_stmt_9250_to_assign_stmt_9254/slice_9249_Update/ca
      -- CP-element group 2: 	 assign_stmt_9250_to_assign_stmt_9254/slice_9253_sample_start_
      -- CP-element group 2: 	 assign_stmt_9250_to_assign_stmt_9254/slice_9253_sample_completed_
      -- CP-element group 2: 	 assign_stmt_9250_to_assign_stmt_9254/slice_9253_update_start_
      -- CP-element group 2: 	 assign_stmt_9250_to_assign_stmt_9254/slice_9253_update_completed_
      -- CP-element group 2: 	 assign_stmt_9250_to_assign_stmt_9254/R_Z_9252_sample_start_
      -- CP-element group 2: 	 assign_stmt_9250_to_assign_stmt_9254/R_Z_9252_sample_completed_
      -- CP-element group 2: 	 assign_stmt_9250_to_assign_stmt_9254/R_Z_9252_update_start_
      -- CP-element group 2: 	 assign_stmt_9250_to_assign_stmt_9254/R_Z_9252_update_completed_
      -- CP-element group 2: 	 assign_stmt_9250_to_assign_stmt_9254/slice_9253_Sample/$entry
      -- CP-element group 2: 	 assign_stmt_9250_to_assign_stmt_9254/slice_9253_Sample/$exit
      -- CP-element group 2: 	 assign_stmt_9250_to_assign_stmt_9254/slice_9253_Sample/rr
      -- CP-element group 2: 	 assign_stmt_9250_to_assign_stmt_9254/slice_9253_Sample/ra
      -- CP-element group 2: 	 assign_stmt_9250_to_assign_stmt_9254/slice_9253_Update/$entry
      -- CP-element group 2: 	 assign_stmt_9250_to_assign_stmt_9254/slice_9253_Update/$exit
      -- CP-element group 2: 	 assign_stmt_9250_to_assign_stmt_9254/slice_9253_Update/cr
      -- CP-element group 2: 	 assign_stmt_9250_to_assign_stmt_9254/slice_9253_Update/ca
      -- CP-element group 2: 	 assign_stmt_9257/$entry
      -- CP-element group 2: 	 assign_stmt_9257/R_Ya_9256_sample_start_
      -- CP-element group 2: 	 assign_stmt_9257/R_Ya_9256_sample_completed_
      -- CP-element group 2: 	 assign_stmt_9257/R_Ya_9256_update_start_
      -- CP-element group 2: 	 assign_stmt_9257/R_Ya_9256_update_completed_
      -- CP-element group 2: 	 assign_stmt_9257/WPIPE_out_data_9255_sample_start_
      -- CP-element group 2: 	 assign_stmt_9257/WPIPE_out_data_9255_Sample/$entry
      -- CP-element group 2: 	 assign_stmt_9257/WPIPE_out_data_9255_Sample/req
      -- 
    -- logger for CP element group c_block_daemon_out_CP_91_elements(2)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and c_block_daemon_out_CP_91_elements(2)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:c_block_daemon_out:CP:c_block_daemon_out_CP_91_elements(2) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:c_block_daemon_out:CP:RPIPE_out_buf_9245_inst_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:c_block_daemon_out:CP:WPIPE_out_data_9255_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ca_110_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_out_buf_9245_inst_ack_1, ack => c_block_daemon_out_CP_91_elements(2)); -- 
    req_164_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => c_block_daemon_out_CP_91_elements(2), ack => WPIPE_out_data_9255_inst_req_0); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 assign_stmt_9257/WPIPE_out_data_9255_sample_completed_
      -- CP-element group 3: 	 assign_stmt_9257/WPIPE_out_data_9255_update_start_
      -- CP-element group 3: 	 assign_stmt_9257/WPIPE_out_data_9255_Sample/$exit
      -- CP-element group 3: 	 assign_stmt_9257/WPIPE_out_data_9255_Sample/ack
      -- CP-element group 3: 	 assign_stmt_9257/WPIPE_out_data_9255_Update/$entry
      -- CP-element group 3: 	 assign_stmt_9257/WPIPE_out_data_9255_Update/req
      -- 
    -- logger for CP element group c_block_daemon_out_CP_91_elements(3)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and c_block_daemon_out_CP_91_elements(3)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:c_block_daemon_out:CP:c_block_daemon_out_CP_91_elements(3) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:c_block_daemon_out:CP:WPIPE_out_data_9255_inst_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:c_block_daemon_out:CP:WPIPE_out_data_9255_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_165_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_out_data_9255_inst_ack_0, ack => c_block_daemon_out_CP_91_elements(3)); -- 
    req_169_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => c_block_daemon_out_CP_91_elements(3), ack => WPIPE_out_data_9255_inst_req_1); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (12) 
      -- CP-element group 4: 	 assign_stmt_9257/$exit
      -- CP-element group 4: 	 assign_stmt_9257/WPIPE_out_data_9255_update_completed_
      -- CP-element group 4: 	 assign_stmt_9257/WPIPE_out_data_9255_Update/$exit
      -- CP-element group 4: 	 assign_stmt_9257/WPIPE_out_data_9255_Update/ack
      -- CP-element group 4: 	 assign_stmt_9260/$entry
      -- CP-element group 4: 	 assign_stmt_9260/R_Yb_9259_sample_start_
      -- CP-element group 4: 	 assign_stmt_9260/R_Yb_9259_sample_completed_
      -- CP-element group 4: 	 assign_stmt_9260/R_Yb_9259_update_start_
      -- CP-element group 4: 	 assign_stmt_9260/R_Yb_9259_update_completed_
      -- CP-element group 4: 	 assign_stmt_9260/WPIPE_out_data_9258_sample_start_
      -- CP-element group 4: 	 assign_stmt_9260/WPIPE_out_data_9258_Sample/$entry
      -- CP-element group 4: 	 assign_stmt_9260/WPIPE_out_data_9258_Sample/req
      -- 
    -- logger for CP element group c_block_daemon_out_CP_91_elements(4)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and c_block_daemon_out_CP_91_elements(4)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:c_block_daemon_out:CP:c_block_daemon_out_CP_91_elements(4) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:c_block_daemon_out:CP:WPIPE_out_data_9255_inst_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:c_block_daemon_out:CP:WPIPE_out_data_9258_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_170_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_out_data_9255_inst_ack_1, ack => c_block_daemon_out_CP_91_elements(4)); -- 
    req_185_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => c_block_daemon_out_CP_91_elements(4), ack => WPIPE_out_data_9258_inst_req_0); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 assign_stmt_9260/WPIPE_out_data_9258_sample_completed_
      -- CP-element group 5: 	 assign_stmt_9260/WPIPE_out_data_9258_update_start_
      -- CP-element group 5: 	 assign_stmt_9260/WPIPE_out_data_9258_Sample/$exit
      -- CP-element group 5: 	 assign_stmt_9260/WPIPE_out_data_9258_Sample/ack
      -- CP-element group 5: 	 assign_stmt_9260/WPIPE_out_data_9258_Update/$entry
      -- CP-element group 5: 	 assign_stmt_9260/WPIPE_out_data_9258_Update/req
      -- 
    -- logger for CP element group c_block_daemon_out_CP_91_elements(5)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and c_block_daemon_out_CP_91_elements(5)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:c_block_daemon_out:CP:c_block_daemon_out_CP_91_elements(5) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:c_block_daemon_out:CP:WPIPE_out_data_9258_inst_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:c_block_daemon_out:CP:WPIPE_out_data_9258_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_186_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_out_data_9258_inst_ack_0, ack => c_block_daemon_out_CP_91_elements(5)); -- 
    req_190_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => c_block_daemon_out_CP_91_elements(5), ack => WPIPE_out_data_9258_inst_req_1); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (5) 
      -- CP-element group 6: 	 $exit
      -- CP-element group 6: 	 assign_stmt_9260/$exit
      -- CP-element group 6: 	 assign_stmt_9260/WPIPE_out_data_9258_update_completed_
      -- CP-element group 6: 	 assign_stmt_9260/WPIPE_out_data_9258_Update/$exit
      -- CP-element group 6: 	 assign_stmt_9260/WPIPE_out_data_9258_Update/ack
      -- 
    -- logger for CP element group c_block_daemon_out_CP_91_elements(6)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and c_block_daemon_out_CP_91_elements(6)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:c_block_daemon_out:CP:c_block_daemon_out_CP_91_elements(6) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:c_block_daemon_out:CP:WPIPE_out_data_9258_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_191_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_out_data_9258_inst_ack_1, ack => c_block_daemon_out_CP_91_elements(6)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal Ya_9250 : std_logic_vector(63 downto 0);
    signal Yb_9254 : std_logic_vector(63 downto 0);
    signal Z_9246 : std_logic_vector(127 downto 0);
    -- 
  begin -- 
    -- logger for split-operator slice_9249_inst flow-through 
    process(Ya_9250) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:c_block_daemon_out:DP:slice_9249_inst:flowthrough inputs: " & " Z_9246 = "& Convert_SLV_To_Hex_String(Z_9246) & " outputs:" & " Ya_9250= "  & Convert_SLV_To_Hex_String(Ya_9250));
      --
    end process; 
    -- flow-through slice operator slice_9249_inst
    Ya_9250 <= Z_9246(127 downto 64);
    -- logger for split-operator slice_9253_inst flow-through 
    process(Yb_9254) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:c_block_daemon_out:DP:slice_9253_inst:flowthrough inputs: " & " Z_9246 = "& Convert_SLV_To_Hex_String(Z_9246) & " outputs:" & " Yb_9254= "  & Convert_SLV_To_Hex_String(Yb_9254));
      --
    end process; 
    -- flow-through slice operator slice_9253_inst
    Yb_9254 <= Z_9246(63 downto 0);
    -- logger for split-operator RPIPE_out_buf_9245_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if RPIPE_out_buf_9245_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:c_block_daemon_out:DP:RPIPE_out_buf_9245_inst:started:   PipeRead from out_buf inputs: " & " no-guard, no-inputs ");
          --
        end if; 
        if RPIPE_out_buf_9245_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:c_block_daemon_out:DP:RPIPE_out_buf_9245_inst:finished:  outputs: " & " Z_9246= "  & Convert_SLV_To_Hex_String(Z_9246));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared inport operator group (0) : RPIPE_out_buf_9245_inst 
    InportGroup0: Block -- 
      signal data_out: std_logic_vector(127 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_out_buf_9245_inst_req_0;
      RPIPE_out_buf_9245_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_out_buf_9245_inst_req_1;
      RPIPE_out_buf_9245_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Z_9246 <= data_out(127 downto 0);
      out_buf_read_0: InputPortRevised -- 
        generic map ( name => "out_buf_read_0", data_width => 128,  num_reqs => 1,  output_buffering => outBUFs,   no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => out_buf_pipe_read_req(0),
          oack => out_buf_pipe_read_ack(0),
          odata => out_buf_pipe_read_data(127 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- logger for split-operator WPIPE_out_data_9255_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if WPIPE_out_data_9255_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:c_block_daemon_out:DP:WPIPE_out_data_9255_inst:started:   PipeWrite to out_data inputs: " & " Ya_9250 = "& Convert_SLV_To_Hex_String(Ya_9250));
          --
        end if; 
        if WPIPE_out_data_9255_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:c_block_daemon_out:DP:WPIPE_out_data_9255_inst:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator WPIPE_out_data_9258_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if WPIPE_out_data_9258_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:c_block_daemon_out:DP:WPIPE_out_data_9258_inst:started:   PipeWrite to out_data inputs: " & " Yb_9254 = "& Convert_SLV_To_Hex_String(Yb_9254));
          --
        end if; 
        if WPIPE_out_data_9258_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:c_block_daemon_out:DP:WPIPE_out_data_9258_inst:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared outport operator group (0) : WPIPE_out_data_9255_inst WPIPE_out_data_9258_inst 
    OutportGroup0: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal sample_req, sample_ack : BooleanArray( 1 downto 0);
      signal update_req, update_ack : BooleanArray( 1 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 1 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      sample_req_unguarded(1) <= WPIPE_out_data_9255_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_out_data_9258_inst_req_0;
      WPIPE_out_data_9255_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_out_data_9258_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(1) <= WPIPE_out_data_9255_inst_req_1;
      update_req_unguarded(0) <= WPIPE_out_data_9258_inst_req_1;
      WPIPE_out_data_9255_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_out_data_9258_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      gI: SplitGuardInterface generic map(nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      data_in <= Ya_9250 & Yb_9254;
      out_data_write_0: OutputPortRevised -- 
        generic map ( name => "out_data", data_width => 64, num_reqs => 2, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => out_data_pipe_write_req(0),
          oack => out_data_pipe_write_ack(0),
          odata => out_data_pipe_write_data(63 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end c_block_daemon_out_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library GhdlLink;
use GhdlLink.LogUtilities.all;
library work;
use work.ahir_system_global_package.all;
entity d_block_daemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    in_buf_pipe_read_req : out  std_logic_vector(0 downto 0);
    in_buf_pipe_read_ack : in   std_logic_vector(0 downto 0);
    in_buf_pipe_read_data : in   std_logic_vector(127 downto 0);
    out_buf_pipe_write_req : out  std_logic_vector(0 downto 0);
    out_buf_pipe_write_ack : in   std_logic_vector(0 downto 0);
    out_buf_pipe_write_data : out  std_logic_vector(127 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity d_block_daemon;
architecture d_block_daemon_arch of d_block_daemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal d_block_daemon_CP_3326_start: Boolean;
  signal d_block_daemon_CP_3326_symbol: Boolean;
  -- volatile/operator module components. 
  component dec_round_Operator is -- 
    port ( -- 
      sample_req: in boolean;
      sample_ack: out boolean;
      update_req: in boolean;
      update_ack: out boolean;
      round_in : in  std_logic_vector(127 downto 0);
      key_in : in  std_logic_vector(127 downto 0);
      l_round : in  std_logic_vector(0 downto 0);
      round_out : out  std_logic_vector(127 downto 0);
      clk, reset: in std_logic
      -- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal W_round_S10_9984_delayed_1_9984_inst_req_1 : boolean;
  signal call_stmt_9991_call_req_0 : boolean;
  signal call_stmt_9991_call_ack_0 : boolean;
  signal call_stmt_9996_call_req_0 : boolean;
  signal W_round_S10_9984_delayed_1_9984_inst_req_0 : boolean;
  signal call_stmt_9991_call_req_1 : boolean;
  signal W_round_S10_9984_delayed_1_9984_inst_ack_0 : boolean;
  signal W_round_S10_9984_delayed_1_9984_inst_ack_1 : boolean;
  signal call_stmt_9991_call_ack_1 : boolean;
  signal call_stmt_9996_call_ack_0 : boolean;
  signal call_stmt_9996_call_req_1 : boolean;
  signal call_stmt_9996_call_ack_1 : boolean;
  signal do_while_stmt_9974_branch_req_0 : boolean;
  signal RPIPE_in_buf_9977_inst_req_0 : boolean;
  signal RPIPE_in_buf_9977_inst_ack_0 : boolean;
  signal RPIPE_in_buf_9977_inst_req_1 : boolean;
  signal RPIPE_in_buf_9977_inst_ack_1 : boolean;
  signal call_stmt_10001_call_req_0 : boolean;
  signal call_stmt_10001_call_ack_0 : boolean;
  signal call_stmt_10001_call_req_1 : boolean;
  signal call_stmt_10001_call_ack_1 : boolean;
  signal call_stmt_10006_call_req_0 : boolean;
  signal call_stmt_10006_call_ack_0 : boolean;
  signal call_stmt_10006_call_req_1 : boolean;
  signal call_stmt_10006_call_ack_1 : boolean;
  signal call_stmt_10011_call_req_0 : boolean;
  signal call_stmt_10011_call_ack_0 : boolean;
  signal call_stmt_10011_call_req_1 : boolean;
  signal call_stmt_10011_call_ack_1 : boolean;
  signal call_stmt_10016_call_req_0 : boolean;
  signal call_stmt_10016_call_ack_0 : boolean;
  signal call_stmt_10016_call_req_1 : boolean;
  signal call_stmt_10016_call_ack_1 : boolean;
  signal call_stmt_10021_call_req_0 : boolean;
  signal call_stmt_10021_call_ack_0 : boolean;
  signal call_stmt_10021_call_req_1 : boolean;
  signal call_stmt_10021_call_ack_1 : boolean;
  signal call_stmt_10026_call_req_0 : boolean;
  signal call_stmt_10026_call_ack_0 : boolean;
  signal call_stmt_10026_call_req_1 : boolean;
  signal call_stmt_10026_call_ack_1 : boolean;
  signal call_stmt_10031_call_req_0 : boolean;
  signal call_stmt_10031_call_ack_0 : boolean;
  signal call_stmt_10031_call_req_1 : boolean;
  signal call_stmt_10031_call_ack_1 : boolean;
  signal call_stmt_10036_call_req_0 : boolean;
  signal call_stmt_10036_call_ack_0 : boolean;
  signal call_stmt_10036_call_req_1 : boolean;
  signal call_stmt_10036_call_ack_1 : boolean;
  signal WPIPE_out_buf_10037_inst_req_0 : boolean;
  signal WPIPE_out_buf_10037_inst_ack_0 : boolean;
  signal WPIPE_out_buf_10037_inst_req_1 : boolean;
  signal WPIPE_out_buf_10037_inst_ack_1 : boolean;
  signal do_while_stmt_9974_branch_ack_0 : boolean;
  signal do_while_stmt_9974_branch_ack_1 : boolean;
  signal global_clock_cycle_count: integer := 0;
  -- 
begin --  
  ---------------------------------------------------------- 
  process(clk)  
  begin -- 
    if(clk'event and clk = '1') then -- 
      if(reset = '1') then -- 
        global_clock_cycle_count <= 0; --
      else -- 
        global_clock_cycle_count <= global_clock_cycle_count + 1; -- 
      end if; --
    end if; --
  end process;
  ---------------------------------------------------------- 
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "d_block_daemon_input_buffer", -- 
      buffer_size => 1,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  d_block_daemon_CP_3326_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "d_block_daemon_out_buffer", -- 
      buffer_size => 1,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= d_block_daemon_CP_3326_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= d_block_daemon_CP_3326_start & tag_ilock_write_ack_symbol;
    gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= d_block_daemon_CP_3326_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  --- logging ------------------------------------------------------
  LogCPEvent(clk,reset,global_clock_cycle_count,d_block_daemon_CP_3326_start,"d_block_daemon cp_entry_symbol ");
  LogCPEvent(clk,reset,global_clock_cycle_count,d_block_daemon_CP_3326_symbol, "d_block_daemon cp_exit_symbol ");
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  d_block_daemon_CP_3326: Block -- control-path 
    signal d_block_daemon_CP_3326_elements: BooleanArray(69 downto 0);
    -- 
  begin -- 
    d_block_daemon_CP_3326_elements(0) <= d_block_daemon_CP_3326_start;
    d_block_daemon_CP_3326_symbol <= d_block_daemon_CP_3326_elements(69);
    -- CP-element group 0:  transition  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (2) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_9973/$entry
      -- 
    -- logger for CP element group d_block_daemon_CP_3326_elements(0)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and d_block_daemon_CP_3326_elements(0)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:d_block_daemon_CP_3326_elements(0) fired."); 
        -- 
      end if; --
    end process; 
    -- CP-element group 1:  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	3 
    -- CP-element group 1:  members (2) 
      -- CP-element group 1: 	 branch_block_stmt_9973/branch_block_stmt_9973__entry__
      -- CP-element group 1: 	 branch_block_stmt_9973/do_while_stmt_9974__entry__
      -- 
    -- logger for CP element group d_block_daemon_CP_3326_elements(1)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and d_block_daemon_CP_3326_elements(1)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:d_block_daemon_CP_3326_elements(1) fired."); 
        -- 
      end if; --
    end process; 
    d_block_daemon_CP_3326_elements(1) <= d_block_daemon_CP_3326_elements(0);
    -- CP-element group 2:  place  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	68 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	69 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_9973/branch_block_stmt_9973__exit__
      -- CP-element group 2: 	 branch_block_stmt_9973/do_while_stmt_9974__exit__
      -- 
    -- logger for CP element group d_block_daemon_CP_3326_elements(2)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and d_block_daemon_CP_3326_elements(2)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:d_block_daemon_CP_3326_elements(2) fired."); 
        -- 
      end if; --
    end process; 
    d_block_daemon_CP_3326_elements(2) <= d_block_daemon_CP_3326_elements(68);
    -- CP-element group 3:  transition  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	1 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_9973/do_while_stmt_9974/$entry
      -- 
    -- logger for CP element group d_block_daemon_CP_3326_elements(3)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and d_block_daemon_CP_3326_elements(3)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:d_block_daemon_CP_3326_elements(3) fired."); 
        -- 
      end if; --
    end process; 
    d_block_daemon_CP_3326_elements(3) <= d_block_daemon_CP_3326_elements(1);
    -- CP-element group 4:  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	10 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974__entry__
      -- 
    -- logger for CP element group d_block_daemon_CP_3326_elements(4)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and d_block_daemon_CP_3326_elements(4)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:d_block_daemon_CP_3326_elements(4) fired."); 
        -- 
      end if; --
    end process; 
    d_block_daemon_CP_3326_elements(4) <= d_block_daemon_CP_3326_elements(3);
    -- CP-element group 5:  merge  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	68 
    -- CP-element group 5:  members (1) 
      -- CP-element group 5: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974__exit__
      -- 
    -- logger for CP element group d_block_daemon_CP_3326_elements(5)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and d_block_daemon_CP_3326_elements(5)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:d_block_daemon_CP_3326_elements(5) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group d_block_daemon_CP_3326_elements(5) is bound as output of CP function.
    -- CP-element group 6:  merge  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	9 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_9973/do_while_stmt_9974/loop_back
      -- 
    -- logger for CP element group d_block_daemon_CP_3326_elements(6)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and d_block_daemon_CP_3326_elements(6)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:d_block_daemon_CP_3326_elements(6) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group d_block_daemon_CP_3326_elements(6) is bound as output of CP function.
    -- CP-element group 7:  branch  place  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	11 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	64 
    -- CP-element group 7: 	66 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_9973/do_while_stmt_9974/condition_done
      -- 
    -- logger for CP element group d_block_daemon_CP_3326_elements(7)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and d_block_daemon_CP_3326_elements(7)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:d_block_daemon_CP_3326_elements(7) fired."); 
        -- 
      end if; --
    end process; 
    d_block_daemon_CP_3326_elements(7) <= d_block_daemon_CP_3326_elements(11);
    -- CP-element group 8:  branch  place  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	63 
    -- CP-element group 8: successors 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_9973/do_while_stmt_9974/loop_body_done
      -- 
    -- logger for CP element group d_block_daemon_CP_3326_elements(8)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and d_block_daemon_CP_3326_elements(8)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:d_block_daemon_CP_3326_elements(8) fired."); 
        -- 
      end if; --
    end process; 
    d_block_daemon_CP_3326_elements(8) <= d_block_daemon_CP_3326_elements(63);
    -- CP-element group 9:  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	6 
    -- CP-element group 9: successors 
    -- CP-element group 9:  members (1) 
      -- CP-element group 9: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/back_edge_to_loop_body
      -- 
    -- logger for CP element group d_block_daemon_CP_3326_elements(9)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and d_block_daemon_CP_3326_elements(9)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:d_block_daemon_CP_3326_elements(9) fired."); 
        -- 
      end if; --
    end process; 
    d_block_daemon_CP_3326_elements(9) <= d_block_daemon_CP_3326_elements(6);
    -- CP-element group 10:  transition  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	4 
    -- CP-element group 10: successors 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/first_time_through_loop_body
      -- 
    -- logger for CP element group d_block_daemon_CP_3326_elements(10)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and d_block_daemon_CP_3326_elements(10)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:d_block_daemon_CP_3326_elements(10) fired."); 
        -- 
      end if; --
    end process; 
    d_block_daemon_CP_3326_elements(10) <= d_block_daemon_CP_3326_elements(4);
    -- CP-element group 11:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	53 
    -- CP-element group 11: 	57 
    -- CP-element group 11: 	7 
    -- CP-element group 11: 	12 
    -- CP-element group 11: 	41 
    -- CP-element group 11: 	45 
    -- CP-element group 11: 	49 
    -- CP-element group 11: 	17 
    -- CP-element group 11: 	21 
    -- CP-element group 11: 	25 
    -- CP-element group 11: 	29 
    -- CP-element group 11: 	33 
    -- CP-element group 11: 	37 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/$entry
      -- CP-element group 11: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/loop_body_start
      -- CP-element group 11: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/condition_evaluated
      -- 
    -- logger for CP element group d_block_daemon_CP_3326_elements(11)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and d_block_daemon_CP_3326_elements(11)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:d_block_daemon_CP_3326_elements(11) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:do_while_stmt_9974_branch_req_0 fired."); 
        -- 
      end if; --
    end process; 
    condition_evaluated_3350_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_3326_elements(11), ack => do_while_stmt_9974_branch_req_0); -- 
    -- Element group d_block_daemon_CP_3326_elements(11) is bound as output of CP function.
    -- CP-element group 12:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: marked-predecessors 
    -- CP-element group 12: 	14 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	14 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/RPIPE_in_buf_9977_sample_start_
      -- CP-element group 12: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/RPIPE_in_buf_9977_Sample/$entry
      -- CP-element group 12: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/RPIPE_in_buf_9977_Sample/rr
      -- 
    -- logger for CP element group d_block_daemon_CP_3326_elements(12)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and d_block_daemon_CP_3326_elements(12)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:d_block_daemon_CP_3326_elements(12) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:RPIPE_in_buf_9977_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_3359_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_3326_elements(12), ack => RPIPE_in_buf_9977_inst_req_0); -- 
    d_block_daemon_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 10,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 34) := "d_block_daemon_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= d_block_daemon_CP_3326_elements(11) & d_block_daemon_CP_3326_elements(14);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => d_block_daemon_CP_3326_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	14 
    -- CP-element group 13: marked-predecessors 
    -- CP-element group 13: 	18 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	15 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/RPIPE_in_buf_9977_update_start_
      -- CP-element group 13: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/RPIPE_in_buf_9977_Update/$entry
      -- CP-element group 13: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/RPIPE_in_buf_9977_Update/cr
      -- 
    -- logger for CP element group d_block_daemon_CP_3326_elements(13)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and d_block_daemon_CP_3326_elements(13)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:d_block_daemon_CP_3326_elements(13) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:RPIPE_in_buf_9977_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_3364_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_3326_elements(13), ack => RPIPE_in_buf_9977_inst_req_1); -- 
    d_block_daemon_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 10,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "d_block_daemon_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= d_block_daemon_CP_3326_elements(14) & d_block_daemon_CP_3326_elements(18);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => d_block_daemon_CP_3326_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	12 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	12 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/RPIPE_in_buf_9977_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/RPIPE_in_buf_9977_Sample/$exit
      -- CP-element group 14: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/RPIPE_in_buf_9977_Sample/ra
      -- 
    -- logger for CP element group d_block_daemon_CP_3326_elements(14)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and d_block_daemon_CP_3326_elements(14)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:d_block_daemon_CP_3326_elements(14) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:RPIPE_in_buf_9977_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_3360_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_in_buf_9977_inst_ack_0, ack => d_block_daemon_CP_3326_elements(14)); -- 
    -- CP-element group 15:  transition  input  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	13 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (23) 
      -- CP-element group 15: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/RPIPE_in_buf_9977_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/RPIPE_in_buf_9977_Update/$exit
      -- CP-element group 15: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/RPIPE_in_buf_9977_Update/ca
      -- CP-element group 15: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/XOR_u128_u128_9982_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/XOR_u128_u128_9982_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/XOR_u128_u128_9982_update_start_
      -- CP-element group 15: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/XOR_u128_u128_9982_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/R_in128_9980_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/R_in128_9980_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/R_in128_9980_update_start_
      -- CP-element group 15: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/R_in128_9980_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/XOR_u128_u128_9982_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/XOR_u128_u128_9982_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/XOR_u128_u128_9982_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/XOR_u128_u128_9982_Sample/ra
      -- CP-element group 15: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/XOR_u128_u128_9982_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/XOR_u128_u128_9982_Update/$exit
      -- CP-element group 15: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/XOR_u128_u128_9982_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/XOR_u128_u128_9982_Update/ca
      -- CP-element group 15: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/R_round_S10_9985_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/R_round_S10_9985_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/R_round_S10_9985_update_start_
      -- CP-element group 15: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/R_round_S10_9985_update_completed_
      -- 
    -- logger for CP element group d_block_daemon_CP_3326_elements(15)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and d_block_daemon_CP_3326_elements(15)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:d_block_daemon_CP_3326_elements(15) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:RPIPE_in_buf_9977_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_3365_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_in_buf_9977_inst_ack_1, ack => d_block_daemon_CP_3326_elements(15)); -- 
    -- CP-element group 16:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	18 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	18 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/assign_stmt_9986_Sample/req
      -- CP-element group 16: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/assign_stmt_9986_sample_start_
      -- CP-element group 16: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/assign_stmt_9986_Sample/$entry
      -- 
    -- logger for CP element group d_block_daemon_CP_3326_elements(16)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and d_block_daemon_CP_3326_elements(16)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:d_block_daemon_CP_3326_elements(16) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:W_round_S10_9984_delayed_1_9984_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_3395_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_3326_elements(16), ack => W_round_S10_9984_delayed_1_9984_inst_req_0); -- 
    d_block_daemon_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 10,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 34) := "d_block_daemon_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= d_block_daemon_CP_3326_elements(15) & d_block_daemon_CP_3326_elements(18);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => d_block_daemon_CP_3326_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	11 
    -- CP-element group 17: marked-predecessors 
    -- CP-element group 17: 	22 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	19 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/assign_stmt_9986_Update/req
      -- CP-element group 17: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/assign_stmt_9986_Update/$entry
      -- CP-element group 17: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/assign_stmt_9986_update_start_
      -- 
    -- logger for CP element group d_block_daemon_CP_3326_elements(17)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and d_block_daemon_CP_3326_elements(17)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:d_block_daemon_CP_3326_elements(17) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:W_round_S10_9984_delayed_1_9984_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_3400_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_3326_elements(17), ack => W_round_S10_9984_delayed_1_9984_inst_req_1); -- 
    d_block_daemon_cp_element_group_17: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 10,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "d_block_daemon_cp_element_group_17"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= d_block_daemon_CP_3326_elements(11) & d_block_daemon_CP_3326_elements(22);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => d_block_daemon_CP_3326_elements(17), clk => clk, reset => reset); --
    end block;
    -- CP-element group 18:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	16 
    -- CP-element group 18: successors 
    -- CP-element group 18: marked-successors 
    -- CP-element group 18: 	13 
    -- CP-element group 18: 	16 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/assign_stmt_9986_Sample/$exit
      -- CP-element group 18: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/assign_stmt_9986_Sample/ack
      -- CP-element group 18: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/assign_stmt_9986_sample_completed_
      -- 
    -- logger for CP element group d_block_daemon_CP_3326_elements(18)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and d_block_daemon_CP_3326_elements(18)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:d_block_daemon_CP_3326_elements(18) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:W_round_S10_9984_delayed_1_9984_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_3396_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => W_round_S10_9984_delayed_1_9984_inst_ack_0, ack => d_block_daemon_CP_3326_elements(18)); -- 
    -- CP-element group 19:  transition  input  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	17 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19:  members (7) 
      -- CP-element group 19: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/assign_stmt_9986_Update/$exit
      -- CP-element group 19: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/R_round_S10_9984_delayed_1_9987_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/R_round_S10_9984_delayed_1_9987_update_start_
      -- CP-element group 19: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/R_round_S10_9984_delayed_1_9987_update_completed_
      -- CP-element group 19: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/R_round_S10_9984_delayed_1_9987_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/assign_stmt_9986_Update/ack
      -- CP-element group 19: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/assign_stmt_9986_update_completed_
      -- 
    -- logger for CP element group d_block_daemon_CP_3326_elements(19)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and d_block_daemon_CP_3326_elements(19)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:d_block_daemon_CP_3326_elements(19) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:W_round_S10_9984_delayed_1_9984_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_3401_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => W_round_S10_9984_delayed_1_9984_inst_ack_1, ack => d_block_daemon_CP_3326_elements(19)); -- 
    -- CP-element group 20:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: marked-predecessors 
    -- CP-element group 20: 	22 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	22 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_9991_Sample/$entry
      -- CP-element group 20: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_9991_Sample/crr
      -- CP-element group 20: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_9991_sample_start_
      -- 
    -- logger for CP element group d_block_daemon_CP_3326_elements(20)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and d_block_daemon_CP_3326_elements(20)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:d_block_daemon_CP_3326_elements(20) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:call_stmt_9991_call_req_0 fired."); 
        -- 
      end if; --
    end process; 
    crr_3413_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_3326_elements(20), ack => call_stmt_9991_call_req_0); -- 
    d_block_daemon_cp_element_group_20: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 10,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 34) := "d_block_daemon_cp_element_group_20"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= d_block_daemon_CP_3326_elements(19) & d_block_daemon_CP_3326_elements(22);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => d_block_daemon_CP_3326_elements(20), clk => clk, reset => reset); --
    end block;
    -- CP-element group 21:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	11 
    -- CP-element group 21: marked-predecessors 
    -- CP-element group 21: 	26 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	23 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_9991_update_start_
      -- CP-element group 21: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_9991_Update/$entry
      -- CP-element group 21: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_9991_Update/ccr
      -- 
    -- logger for CP element group d_block_daemon_CP_3326_elements(21)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and d_block_daemon_CP_3326_elements(21)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:d_block_daemon_CP_3326_elements(21) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:call_stmt_9991_call_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ccr_3418_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_3326_elements(21), ack => call_stmt_9991_call_req_1); -- 
    d_block_daemon_cp_element_group_21: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 10,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "d_block_daemon_cp_element_group_21"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= d_block_daemon_CP_3326_elements(11) & d_block_daemon_CP_3326_elements(26);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => d_block_daemon_CP_3326_elements(21), clk => clk, reset => reset); --
    end block;
    -- CP-element group 22:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	20 
    -- CP-element group 22: successors 
    -- CP-element group 22: marked-successors 
    -- CP-element group 22: 	17 
    -- CP-element group 22: 	20 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_9991_Sample/$exit
      -- CP-element group 22: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_9991_Sample/cra
      -- CP-element group 22: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_9991_sample_completed_
      -- 
    -- logger for CP element group d_block_daemon_CP_3326_elements(22)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and d_block_daemon_CP_3326_elements(22)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:d_block_daemon_CP_3326_elements(22) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:call_stmt_9991_call_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    cra_3414_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_9991_call_ack_0, ack => d_block_daemon_CP_3326_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	21 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	24 
    -- CP-element group 23:  members (7) 
      -- CP-element group 23: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/R_round_S9_9992_sample_completed_
      -- CP-element group 23: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_9991_update_completed_
      -- CP-element group 23: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_9991_Update/$exit
      -- CP-element group 23: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/R_round_S9_9992_update_completed_
      -- CP-element group 23: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/R_round_S9_9992_update_start_
      -- CP-element group 23: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/R_round_S9_9992_sample_start_
      -- CP-element group 23: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_9991_Update/cca
      -- 
    -- logger for CP element group d_block_daemon_CP_3326_elements(23)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and d_block_daemon_CP_3326_elements(23)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:d_block_daemon_CP_3326_elements(23) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:call_stmt_9991_call_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    cca_3419_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_9991_call_ack_1, ack => d_block_daemon_CP_3326_elements(23)); -- 
    -- CP-element group 24:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	23 
    -- CP-element group 24: marked-predecessors 
    -- CP-element group 24: 	26 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	26 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_9996_Sample/$entry
      -- CP-element group 24: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_9996_Sample/crr
      -- CP-element group 24: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_9996_sample_start_
      -- 
    -- logger for CP element group d_block_daemon_CP_3326_elements(24)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and d_block_daemon_CP_3326_elements(24)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:d_block_daemon_CP_3326_elements(24) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:call_stmt_9996_call_req_0 fired."); 
        -- 
      end if; --
    end process; 
    crr_3431_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_3326_elements(24), ack => call_stmt_9996_call_req_0); -- 
    d_block_daemon_cp_element_group_24: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 10,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 34) := "d_block_daemon_cp_element_group_24"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= d_block_daemon_CP_3326_elements(23) & d_block_daemon_CP_3326_elements(26);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => d_block_daemon_CP_3326_elements(24), clk => clk, reset => reset); --
    end block;
    -- CP-element group 25:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	11 
    -- CP-element group 25: marked-predecessors 
    -- CP-element group 25: 	30 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	27 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_9996_update_start_
      -- CP-element group 25: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_9996_Update/$entry
      -- CP-element group 25: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_9996_Update/ccr
      -- 
    -- logger for CP element group d_block_daemon_CP_3326_elements(25)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and d_block_daemon_CP_3326_elements(25)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:d_block_daemon_CP_3326_elements(25) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:call_stmt_9996_call_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ccr_3436_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_3326_elements(25), ack => call_stmt_9996_call_req_1); -- 
    d_block_daemon_cp_element_group_25: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 10,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "d_block_daemon_cp_element_group_25"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= d_block_daemon_CP_3326_elements(11) & d_block_daemon_CP_3326_elements(30);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => d_block_daemon_CP_3326_elements(25), clk => clk, reset => reset); --
    end block;
    -- CP-element group 26:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	24 
    -- CP-element group 26: successors 
    -- CP-element group 26: marked-successors 
    -- CP-element group 26: 	21 
    -- CP-element group 26: 	24 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_9996_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_9996_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_9996_Sample/cra
      -- 
    -- logger for CP element group d_block_daemon_CP_3326_elements(26)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and d_block_daemon_CP_3326_elements(26)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:d_block_daemon_CP_3326_elements(26) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:call_stmt_9996_call_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    cra_3432_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_9996_call_ack_0, ack => d_block_daemon_CP_3326_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	25 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	28 
    -- CP-element group 27:  members (7) 
      -- CP-element group 27: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/R_round_S8_9997_sample_start_
      -- CP-element group 27: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/R_round_S8_9997_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/R_round_S8_9997_update_start_
      -- CP-element group 27: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/R_round_S8_9997_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_9996_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_9996_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_9996_Update/cca
      -- 
    -- logger for CP element group d_block_daemon_CP_3326_elements(27)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and d_block_daemon_CP_3326_elements(27)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:d_block_daemon_CP_3326_elements(27) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:call_stmt_9996_call_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    cca_3437_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_9996_call_ack_1, ack => d_block_daemon_CP_3326_elements(27)); -- 
    -- CP-element group 28:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	27 
    -- CP-element group 28: marked-predecessors 
    -- CP-element group 28: 	30 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	30 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_10001_sample_start_
      -- CP-element group 28: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_10001_Sample/$entry
      -- CP-element group 28: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_10001_Sample/crr
      -- 
    -- logger for CP element group d_block_daemon_CP_3326_elements(28)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and d_block_daemon_CP_3326_elements(28)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:d_block_daemon_CP_3326_elements(28) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:call_stmt_10001_call_req_0 fired."); 
        -- 
      end if; --
    end process; 
    crr_3449_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_3326_elements(28), ack => call_stmt_10001_call_req_0); -- 
    d_block_daemon_cp_element_group_28: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 10,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 34) := "d_block_daemon_cp_element_group_28"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= d_block_daemon_CP_3326_elements(27) & d_block_daemon_CP_3326_elements(30);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => d_block_daemon_CP_3326_elements(28), clk => clk, reset => reset); --
    end block;
    -- CP-element group 29:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	11 
    -- CP-element group 29: marked-predecessors 
    -- CP-element group 29: 	34 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	31 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_10001_update_start_
      -- CP-element group 29: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_10001_Update/$entry
      -- CP-element group 29: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_10001_Update/ccr
      -- 
    -- logger for CP element group d_block_daemon_CP_3326_elements(29)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and d_block_daemon_CP_3326_elements(29)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:d_block_daemon_CP_3326_elements(29) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:call_stmt_10001_call_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ccr_3454_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_3326_elements(29), ack => call_stmt_10001_call_req_1); -- 
    d_block_daemon_cp_element_group_29: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 10,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "d_block_daemon_cp_element_group_29"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= d_block_daemon_CP_3326_elements(11) & d_block_daemon_CP_3326_elements(34);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => d_block_daemon_CP_3326_elements(29), clk => clk, reset => reset); --
    end block;
    -- CP-element group 30:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	28 
    -- CP-element group 30: successors 
    -- CP-element group 30: marked-successors 
    -- CP-element group 30: 	25 
    -- CP-element group 30: 	28 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_10001_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_10001_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_10001_Sample/cra
      -- 
    -- logger for CP element group d_block_daemon_CP_3326_elements(30)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and d_block_daemon_CP_3326_elements(30)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:d_block_daemon_CP_3326_elements(30) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:call_stmt_10001_call_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    cra_3450_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_10001_call_ack_0, ack => d_block_daemon_CP_3326_elements(30)); -- 
    -- CP-element group 31:  transition  input  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	29 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31:  members (7) 
      -- CP-element group 31: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/R_round_S7_10002_sample_completed_
      -- CP-element group 31: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_10001_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_10001_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_10001_Update/cca
      -- CP-element group 31: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/R_round_S7_10002_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/R_round_S7_10002_update_start_
      -- CP-element group 31: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/R_round_S7_10002_update_completed_
      -- 
    -- logger for CP element group d_block_daemon_CP_3326_elements(31)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and d_block_daemon_CP_3326_elements(31)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:d_block_daemon_CP_3326_elements(31) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:call_stmt_10001_call_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    cca_3455_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_10001_call_ack_1, ack => d_block_daemon_CP_3326_elements(31)); -- 
    -- CP-element group 32:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	31 
    -- CP-element group 32: marked-predecessors 
    -- CP-element group 32: 	34 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	34 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_10006_sample_start_
      -- CP-element group 32: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_10006_Sample/$entry
      -- CP-element group 32: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_10006_Sample/crr
      -- 
    -- logger for CP element group d_block_daemon_CP_3326_elements(32)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and d_block_daemon_CP_3326_elements(32)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:d_block_daemon_CP_3326_elements(32) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:call_stmt_10006_call_req_0 fired."); 
        -- 
      end if; --
    end process; 
    crr_3467_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_3326_elements(32), ack => call_stmt_10006_call_req_0); -- 
    d_block_daemon_cp_element_group_32: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 10,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 34) := "d_block_daemon_cp_element_group_32"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= d_block_daemon_CP_3326_elements(31) & d_block_daemon_CP_3326_elements(34);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => d_block_daemon_CP_3326_elements(32), clk => clk, reset => reset); --
    end block;
    -- CP-element group 33:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	11 
    -- CP-element group 33: marked-predecessors 
    -- CP-element group 33: 	38 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	35 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_10006_update_start_
      -- CP-element group 33: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_10006_Update/$entry
      -- CP-element group 33: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_10006_Update/ccr
      -- 
    -- logger for CP element group d_block_daemon_CP_3326_elements(33)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and d_block_daemon_CP_3326_elements(33)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:d_block_daemon_CP_3326_elements(33) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:call_stmt_10006_call_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ccr_3472_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_3326_elements(33), ack => call_stmt_10006_call_req_1); -- 
    d_block_daemon_cp_element_group_33: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 10,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "d_block_daemon_cp_element_group_33"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= d_block_daemon_CP_3326_elements(11) & d_block_daemon_CP_3326_elements(38);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => d_block_daemon_CP_3326_elements(33), clk => clk, reset => reset); --
    end block;
    -- CP-element group 34:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	32 
    -- CP-element group 34: successors 
    -- CP-element group 34: marked-successors 
    -- CP-element group 34: 	29 
    -- CP-element group 34: 	32 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_10006_sample_completed_
      -- CP-element group 34: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_10006_Sample/$exit
      -- CP-element group 34: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_10006_Sample/cra
      -- 
    -- logger for CP element group d_block_daemon_CP_3326_elements(34)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and d_block_daemon_CP_3326_elements(34)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:d_block_daemon_CP_3326_elements(34) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:call_stmt_10006_call_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    cra_3468_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_10006_call_ack_0, ack => d_block_daemon_CP_3326_elements(34)); -- 
    -- CP-element group 35:  transition  input  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	33 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	36 
    -- CP-element group 35:  members (7) 
      -- CP-element group 35: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_10006_update_completed_
      -- CP-element group 35: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_10006_Update/$exit
      -- CP-element group 35: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_10006_Update/cca
      -- CP-element group 35: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/R_round_S6_10007_sample_start_
      -- CP-element group 35: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/R_round_S6_10007_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/R_round_S6_10007_update_start_
      -- CP-element group 35: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/R_round_S6_10007_update_completed_
      -- 
    -- logger for CP element group d_block_daemon_CP_3326_elements(35)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and d_block_daemon_CP_3326_elements(35)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:d_block_daemon_CP_3326_elements(35) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:call_stmt_10006_call_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    cca_3473_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_10006_call_ack_1, ack => d_block_daemon_CP_3326_elements(35)); -- 
    -- CP-element group 36:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	35 
    -- CP-element group 36: marked-predecessors 
    -- CP-element group 36: 	38 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	38 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_10011_sample_start_
      -- CP-element group 36: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_10011_Sample/$entry
      -- CP-element group 36: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_10011_Sample/crr
      -- 
    -- logger for CP element group d_block_daemon_CP_3326_elements(36)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and d_block_daemon_CP_3326_elements(36)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:d_block_daemon_CP_3326_elements(36) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:call_stmt_10011_call_req_0 fired."); 
        -- 
      end if; --
    end process; 
    crr_3485_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_3326_elements(36), ack => call_stmt_10011_call_req_0); -- 
    d_block_daemon_cp_element_group_36: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 10,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 34) := "d_block_daemon_cp_element_group_36"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= d_block_daemon_CP_3326_elements(35) & d_block_daemon_CP_3326_elements(38);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => d_block_daemon_CP_3326_elements(36), clk => clk, reset => reset); --
    end block;
    -- CP-element group 37:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	11 
    -- CP-element group 37: marked-predecessors 
    -- CP-element group 37: 	42 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	39 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_10011_update_start_
      -- CP-element group 37: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_10011_Update/$entry
      -- CP-element group 37: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_10011_Update/ccr
      -- 
    -- logger for CP element group d_block_daemon_CP_3326_elements(37)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and d_block_daemon_CP_3326_elements(37)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:d_block_daemon_CP_3326_elements(37) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:call_stmt_10011_call_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ccr_3490_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_3326_elements(37), ack => call_stmt_10011_call_req_1); -- 
    d_block_daemon_cp_element_group_37: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 10,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "d_block_daemon_cp_element_group_37"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= d_block_daemon_CP_3326_elements(11) & d_block_daemon_CP_3326_elements(42);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => d_block_daemon_CP_3326_elements(37), clk => clk, reset => reset); --
    end block;
    -- CP-element group 38:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	36 
    -- CP-element group 38: successors 
    -- CP-element group 38: marked-successors 
    -- CP-element group 38: 	33 
    -- CP-element group 38: 	36 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_10011_sample_completed_
      -- CP-element group 38: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_10011_Sample/$exit
      -- CP-element group 38: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_10011_Sample/cra
      -- 
    -- logger for CP element group d_block_daemon_CP_3326_elements(38)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and d_block_daemon_CP_3326_elements(38)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:d_block_daemon_CP_3326_elements(38) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:call_stmt_10011_call_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    cra_3486_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_10011_call_ack_0, ack => d_block_daemon_CP_3326_elements(38)); -- 
    -- CP-element group 39:  transition  input  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	37 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	40 
    -- CP-element group 39:  members (7) 
      -- CP-element group 39: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_10011_update_completed_
      -- CP-element group 39: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_10011_Update/$exit
      -- CP-element group 39: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_10011_Update/cca
      -- CP-element group 39: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/R_round_S5_10012_sample_start_
      -- CP-element group 39: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/R_round_S5_10012_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/R_round_S5_10012_update_start_
      -- CP-element group 39: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/R_round_S5_10012_update_completed_
      -- 
    -- logger for CP element group d_block_daemon_CP_3326_elements(39)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and d_block_daemon_CP_3326_elements(39)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:d_block_daemon_CP_3326_elements(39) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:call_stmt_10011_call_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    cca_3491_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_10011_call_ack_1, ack => d_block_daemon_CP_3326_elements(39)); -- 
    -- CP-element group 40:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	39 
    -- CP-element group 40: marked-predecessors 
    -- CP-element group 40: 	42 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	42 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_10016_sample_start_
      -- CP-element group 40: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_10016_Sample/$entry
      -- CP-element group 40: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_10016_Sample/crr
      -- 
    -- logger for CP element group d_block_daemon_CP_3326_elements(40)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and d_block_daemon_CP_3326_elements(40)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:d_block_daemon_CP_3326_elements(40) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:call_stmt_10016_call_req_0 fired."); 
        -- 
      end if; --
    end process; 
    crr_3503_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_3326_elements(40), ack => call_stmt_10016_call_req_0); -- 
    d_block_daemon_cp_element_group_40: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 10,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 34) := "d_block_daemon_cp_element_group_40"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= d_block_daemon_CP_3326_elements(39) & d_block_daemon_CP_3326_elements(42);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => d_block_daemon_CP_3326_elements(40), clk => clk, reset => reset); --
    end block;
    -- CP-element group 41:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	11 
    -- CP-element group 41: marked-predecessors 
    -- CP-element group 41: 	46 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	43 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_10016_update_start_
      -- CP-element group 41: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_10016_Update/$entry
      -- CP-element group 41: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_10016_Update/ccr
      -- 
    -- logger for CP element group d_block_daemon_CP_3326_elements(41)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and d_block_daemon_CP_3326_elements(41)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:d_block_daemon_CP_3326_elements(41) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:call_stmt_10016_call_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ccr_3508_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_3326_elements(41), ack => call_stmt_10016_call_req_1); -- 
    d_block_daemon_cp_element_group_41: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 10,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "d_block_daemon_cp_element_group_41"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= d_block_daemon_CP_3326_elements(11) & d_block_daemon_CP_3326_elements(46);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => d_block_daemon_CP_3326_elements(41), clk => clk, reset => reset); --
    end block;
    -- CP-element group 42:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	40 
    -- CP-element group 42: successors 
    -- CP-element group 42: marked-successors 
    -- CP-element group 42: 	40 
    -- CP-element group 42: 	37 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_10016_sample_completed_
      -- CP-element group 42: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_10016_Sample/$exit
      -- CP-element group 42: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_10016_Sample/cra
      -- 
    -- logger for CP element group d_block_daemon_CP_3326_elements(42)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and d_block_daemon_CP_3326_elements(42)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:d_block_daemon_CP_3326_elements(42) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:call_stmt_10016_call_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    cra_3504_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_10016_call_ack_0, ack => d_block_daemon_CP_3326_elements(42)); -- 
    -- CP-element group 43:  transition  input  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	41 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	44 
    -- CP-element group 43:  members (7) 
      -- CP-element group 43: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_10016_update_completed_
      -- CP-element group 43: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_10016_Update/$exit
      -- CP-element group 43: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_10016_Update/cca
      -- CP-element group 43: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/R_round_S4_10017_sample_start_
      -- CP-element group 43: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/R_round_S4_10017_sample_completed_
      -- CP-element group 43: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/R_round_S4_10017_update_start_
      -- CP-element group 43: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/R_round_S4_10017_update_completed_
      -- 
    -- logger for CP element group d_block_daemon_CP_3326_elements(43)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and d_block_daemon_CP_3326_elements(43)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:d_block_daemon_CP_3326_elements(43) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:call_stmt_10016_call_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    cca_3509_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_10016_call_ack_1, ack => d_block_daemon_CP_3326_elements(43)); -- 
    -- CP-element group 44:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	43 
    -- CP-element group 44: marked-predecessors 
    -- CP-element group 44: 	46 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	46 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_10021_sample_start_
      -- CP-element group 44: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_10021_Sample/$entry
      -- CP-element group 44: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_10021_Sample/crr
      -- 
    -- logger for CP element group d_block_daemon_CP_3326_elements(44)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and d_block_daemon_CP_3326_elements(44)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:d_block_daemon_CP_3326_elements(44) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:call_stmt_10021_call_req_0 fired."); 
        -- 
      end if; --
    end process; 
    crr_3521_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_3326_elements(44), ack => call_stmt_10021_call_req_0); -- 
    d_block_daemon_cp_element_group_44: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 10,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 34) := "d_block_daemon_cp_element_group_44"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= d_block_daemon_CP_3326_elements(43) & d_block_daemon_CP_3326_elements(46);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => d_block_daemon_CP_3326_elements(44), clk => clk, reset => reset); --
    end block;
    -- CP-element group 45:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	11 
    -- CP-element group 45: marked-predecessors 
    -- CP-element group 45: 	50 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	47 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_10021_update_start_
      -- CP-element group 45: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_10021_Update/$entry
      -- CP-element group 45: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_10021_Update/ccr
      -- 
    -- logger for CP element group d_block_daemon_CP_3326_elements(45)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and d_block_daemon_CP_3326_elements(45)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:d_block_daemon_CP_3326_elements(45) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:call_stmt_10021_call_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ccr_3526_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_3326_elements(45), ack => call_stmt_10021_call_req_1); -- 
    d_block_daemon_cp_element_group_45: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 10,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "d_block_daemon_cp_element_group_45"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= d_block_daemon_CP_3326_elements(11) & d_block_daemon_CP_3326_elements(50);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => d_block_daemon_CP_3326_elements(45), clk => clk, reset => reset); --
    end block;
    -- CP-element group 46:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	44 
    -- CP-element group 46: successors 
    -- CP-element group 46: marked-successors 
    -- CP-element group 46: 	41 
    -- CP-element group 46: 	44 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_10021_sample_completed_
      -- CP-element group 46: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_10021_Sample/$exit
      -- CP-element group 46: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_10021_Sample/cra
      -- 
    -- logger for CP element group d_block_daemon_CP_3326_elements(46)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and d_block_daemon_CP_3326_elements(46)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:d_block_daemon_CP_3326_elements(46) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:call_stmt_10021_call_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    cra_3522_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_10021_call_ack_0, ack => d_block_daemon_CP_3326_elements(46)); -- 
    -- CP-element group 47:  transition  input  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	45 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	48 
    -- CP-element group 47:  members (7) 
      -- CP-element group 47: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_10021_update_completed_
      -- CP-element group 47: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_10021_Update/$exit
      -- CP-element group 47: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_10021_Update/cca
      -- CP-element group 47: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/R_round_S3_10022_sample_start_
      -- CP-element group 47: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/R_round_S3_10022_sample_completed_
      -- CP-element group 47: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/R_round_S3_10022_update_start_
      -- CP-element group 47: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/R_round_S3_10022_update_completed_
      -- 
    -- logger for CP element group d_block_daemon_CP_3326_elements(47)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and d_block_daemon_CP_3326_elements(47)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:d_block_daemon_CP_3326_elements(47) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:call_stmt_10021_call_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    cca_3527_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_10021_call_ack_1, ack => d_block_daemon_CP_3326_elements(47)); -- 
    -- CP-element group 48:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	47 
    -- CP-element group 48: marked-predecessors 
    -- CP-element group 48: 	50 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	50 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_10026_sample_start_
      -- CP-element group 48: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_10026_Sample/$entry
      -- CP-element group 48: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_10026_Sample/crr
      -- 
    -- logger for CP element group d_block_daemon_CP_3326_elements(48)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and d_block_daemon_CP_3326_elements(48)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:d_block_daemon_CP_3326_elements(48) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:call_stmt_10026_call_req_0 fired."); 
        -- 
      end if; --
    end process; 
    crr_3539_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_3326_elements(48), ack => call_stmt_10026_call_req_0); -- 
    d_block_daemon_cp_element_group_48: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 10,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 34) := "d_block_daemon_cp_element_group_48"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= d_block_daemon_CP_3326_elements(47) & d_block_daemon_CP_3326_elements(50);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => d_block_daemon_CP_3326_elements(48), clk => clk, reset => reset); --
    end block;
    -- CP-element group 49:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	11 
    -- CP-element group 49: marked-predecessors 
    -- CP-element group 49: 	54 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	51 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_10026_update_start_
      -- CP-element group 49: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_10026_Update/$entry
      -- CP-element group 49: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_10026_Update/ccr
      -- 
    -- logger for CP element group d_block_daemon_CP_3326_elements(49)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and d_block_daemon_CP_3326_elements(49)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:d_block_daemon_CP_3326_elements(49) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:call_stmt_10026_call_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ccr_3544_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_3326_elements(49), ack => call_stmt_10026_call_req_1); -- 
    d_block_daemon_cp_element_group_49: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 10,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "d_block_daemon_cp_element_group_49"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= d_block_daemon_CP_3326_elements(11) & d_block_daemon_CP_3326_elements(54);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => d_block_daemon_CP_3326_elements(49), clk => clk, reset => reset); --
    end block;
    -- CP-element group 50:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	48 
    -- CP-element group 50: successors 
    -- CP-element group 50: marked-successors 
    -- CP-element group 50: 	45 
    -- CP-element group 50: 	48 
    -- CP-element group 50:  members (3) 
      -- CP-element group 50: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_10026_sample_completed_
      -- CP-element group 50: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_10026_Sample/$exit
      -- CP-element group 50: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_10026_Sample/cra
      -- 
    -- logger for CP element group d_block_daemon_CP_3326_elements(50)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and d_block_daemon_CP_3326_elements(50)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:d_block_daemon_CP_3326_elements(50) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:call_stmt_10026_call_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    cra_3540_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_10026_call_ack_0, ack => d_block_daemon_CP_3326_elements(50)); -- 
    -- CP-element group 51:  transition  input  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	49 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	52 
    -- CP-element group 51:  members (7) 
      -- CP-element group 51: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_10026_update_completed_
      -- CP-element group 51: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_10026_Update/$exit
      -- CP-element group 51: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_10026_Update/cca
      -- CP-element group 51: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/R_round_S2_10027_sample_start_
      -- CP-element group 51: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/R_round_S2_10027_sample_completed_
      -- CP-element group 51: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/R_round_S2_10027_update_start_
      -- CP-element group 51: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/R_round_S2_10027_update_completed_
      -- 
    -- logger for CP element group d_block_daemon_CP_3326_elements(51)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and d_block_daemon_CP_3326_elements(51)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:d_block_daemon_CP_3326_elements(51) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:call_stmt_10026_call_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    cca_3545_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_10026_call_ack_1, ack => d_block_daemon_CP_3326_elements(51)); -- 
    -- CP-element group 52:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	51 
    -- CP-element group 52: marked-predecessors 
    -- CP-element group 52: 	54 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	54 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_10031_sample_start_
      -- CP-element group 52: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_10031_Sample/$entry
      -- CP-element group 52: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_10031_Sample/crr
      -- 
    -- logger for CP element group d_block_daemon_CP_3326_elements(52)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and d_block_daemon_CP_3326_elements(52)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:d_block_daemon_CP_3326_elements(52) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:call_stmt_10031_call_req_0 fired."); 
        -- 
      end if; --
    end process; 
    crr_3557_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_3326_elements(52), ack => call_stmt_10031_call_req_0); -- 
    d_block_daemon_cp_element_group_52: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 10,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 34) := "d_block_daemon_cp_element_group_52"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= d_block_daemon_CP_3326_elements(51) & d_block_daemon_CP_3326_elements(54);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => d_block_daemon_CP_3326_elements(52), clk => clk, reset => reset); --
    end block;
    -- CP-element group 53:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	11 
    -- CP-element group 53: marked-predecessors 
    -- CP-element group 53: 	58 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	55 
    -- CP-element group 53:  members (3) 
      -- CP-element group 53: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_10031_update_start_
      -- CP-element group 53: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_10031_Update/$entry
      -- CP-element group 53: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_10031_Update/ccr
      -- 
    -- logger for CP element group d_block_daemon_CP_3326_elements(53)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and d_block_daemon_CP_3326_elements(53)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:d_block_daemon_CP_3326_elements(53) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:call_stmt_10031_call_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ccr_3562_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_3326_elements(53), ack => call_stmt_10031_call_req_1); -- 
    d_block_daemon_cp_element_group_53: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 10,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "d_block_daemon_cp_element_group_53"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= d_block_daemon_CP_3326_elements(11) & d_block_daemon_CP_3326_elements(58);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => d_block_daemon_CP_3326_elements(53), clk => clk, reset => reset); --
    end block;
    -- CP-element group 54:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	52 
    -- CP-element group 54: successors 
    -- CP-element group 54: marked-successors 
    -- CP-element group 54: 	52 
    -- CP-element group 54: 	49 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_10031_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_10031_Sample/$exit
      -- CP-element group 54: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_10031_Sample/cra
      -- 
    -- logger for CP element group d_block_daemon_CP_3326_elements(54)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and d_block_daemon_CP_3326_elements(54)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:d_block_daemon_CP_3326_elements(54) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:call_stmt_10031_call_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    cra_3558_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_10031_call_ack_0, ack => d_block_daemon_CP_3326_elements(54)); -- 
    -- CP-element group 55:  transition  input  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	53 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55:  members (7) 
      -- CP-element group 55: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_10031_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_10031_Update/$exit
      -- CP-element group 55: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_10031_Update/cca
      -- CP-element group 55: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/R_round_S1_10032_sample_start_
      -- CP-element group 55: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/R_round_S1_10032_sample_completed_
      -- CP-element group 55: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/R_round_S1_10032_update_start_
      -- CP-element group 55: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/R_round_S1_10032_update_completed_
      -- 
    -- logger for CP element group d_block_daemon_CP_3326_elements(55)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and d_block_daemon_CP_3326_elements(55)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:d_block_daemon_CP_3326_elements(55) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:call_stmt_10031_call_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    cca_3563_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_10031_call_ack_1, ack => d_block_daemon_CP_3326_elements(55)); -- 
    -- CP-element group 56:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	55 
    -- CP-element group 56: marked-predecessors 
    -- CP-element group 56: 	58 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	58 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_10036_sample_start_
      -- CP-element group 56: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_10036_Sample/$entry
      -- CP-element group 56: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_10036_Sample/crr
      -- 
    -- logger for CP element group d_block_daemon_CP_3326_elements(56)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and d_block_daemon_CP_3326_elements(56)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:d_block_daemon_CP_3326_elements(56) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:call_stmt_10036_call_req_0 fired."); 
        -- 
      end if; --
    end process; 
    crr_3575_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_3326_elements(56), ack => call_stmt_10036_call_req_0); -- 
    d_block_daemon_cp_element_group_56: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 10,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 34) := "d_block_daemon_cp_element_group_56"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= d_block_daemon_CP_3326_elements(55) & d_block_daemon_CP_3326_elements(58);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => d_block_daemon_CP_3326_elements(56), clk => clk, reset => reset); --
    end block;
    -- CP-element group 57:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	11 
    -- CP-element group 57: marked-predecessors 
    -- CP-element group 57: 	62 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	59 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_10036_Update/$entry
      -- CP-element group 57: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_10036_update_start_
      -- CP-element group 57: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_10036_Update/ccr
      -- 
    -- logger for CP element group d_block_daemon_CP_3326_elements(57)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and d_block_daemon_CP_3326_elements(57)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:d_block_daemon_CP_3326_elements(57) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:call_stmt_10036_call_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ccr_3580_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_3326_elements(57), ack => call_stmt_10036_call_req_1); -- 
    d_block_daemon_cp_element_group_57: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 10,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "d_block_daemon_cp_element_group_57"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= d_block_daemon_CP_3326_elements(11) & d_block_daemon_CP_3326_elements(62);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => d_block_daemon_CP_3326_elements(57), clk => clk, reset => reset); --
    end block;
    -- CP-element group 58:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	56 
    -- CP-element group 58: successors 
    -- CP-element group 58: marked-successors 
    -- CP-element group 58: 	53 
    -- CP-element group 58: 	56 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_10036_sample_completed_
      -- CP-element group 58: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_10036_Sample/$exit
      -- CP-element group 58: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_10036_Sample/cra
      -- 
    -- logger for CP element group d_block_daemon_CP_3326_elements(58)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and d_block_daemon_CP_3326_elements(58)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:d_block_daemon_CP_3326_elements(58) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:call_stmt_10036_call_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    cra_3576_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_10036_call_ack_0, ack => d_block_daemon_CP_3326_elements(58)); -- 
    -- CP-element group 59:  transition  input  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	57 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	60 
    -- CP-element group 59:  members (7) 
      -- CP-element group 59: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_10036_update_completed_
      -- CP-element group 59: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_10036_Update/$exit
      -- CP-element group 59: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/call_stmt_10036_Update/cca
      -- CP-element group 59: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/R_round_S0_10038_sample_start_
      -- CP-element group 59: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/R_round_S0_10038_sample_completed_
      -- CP-element group 59: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/R_round_S0_10038_update_start_
      -- CP-element group 59: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/R_round_S0_10038_update_completed_
      -- 
    -- logger for CP element group d_block_daemon_CP_3326_elements(59)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and d_block_daemon_CP_3326_elements(59)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:d_block_daemon_CP_3326_elements(59) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:call_stmt_10036_call_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    cca_3581_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_10036_call_ack_1, ack => d_block_daemon_CP_3326_elements(59)); -- 
    -- CP-element group 60:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	59 
    -- CP-element group 60: marked-predecessors 
    -- CP-element group 60: 	62 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	62 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/WPIPE_out_buf_10037_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/WPIPE_out_buf_10037_Sample/$entry
      -- CP-element group 60: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/WPIPE_out_buf_10037_Sample/req
      -- 
    -- logger for CP element group d_block_daemon_CP_3326_elements(60)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and d_block_daemon_CP_3326_elements(60)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:d_block_daemon_CP_3326_elements(60) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:WPIPE_out_buf_10037_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_3593_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_3326_elements(60), ack => WPIPE_out_buf_10037_inst_req_0); -- 
    d_block_daemon_cp_element_group_60: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 10,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 34) := "d_block_daemon_cp_element_group_60"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= d_block_daemon_CP_3326_elements(59) & d_block_daemon_CP_3326_elements(62);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => d_block_daemon_CP_3326_elements(60), clk => clk, reset => reset); --
    end block;
    -- CP-element group 61:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	62 
    -- CP-element group 61: marked-predecessors 
    -- CP-element group 61: 	63 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	63 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/WPIPE_out_buf_10037_update_start_
      -- CP-element group 61: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/WPIPE_out_buf_10037_Update/$entry
      -- CP-element group 61: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/WPIPE_out_buf_10037_Update/req
      -- 
    -- logger for CP element group d_block_daemon_CP_3326_elements(61)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and d_block_daemon_CP_3326_elements(61)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:d_block_daemon_CP_3326_elements(61) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:WPIPE_out_buf_10037_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_3598_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_3326_elements(61), ack => WPIPE_out_buf_10037_inst_req_1); -- 
    d_block_daemon_cp_element_group_61: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 10,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "d_block_daemon_cp_element_group_61"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= d_block_daemon_CP_3326_elements(62) & d_block_daemon_CP_3326_elements(63);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => d_block_daemon_CP_3326_elements(61), clk => clk, reset => reset); --
    end block;
    -- CP-element group 62:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	60 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	61 
    -- CP-element group 62: marked-successors 
    -- CP-element group 62: 	57 
    -- CP-element group 62: 	60 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/WPIPE_out_buf_10037_sample_completed_
      -- CP-element group 62: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/WPIPE_out_buf_10037_Sample/$exit
      -- CP-element group 62: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/WPIPE_out_buf_10037_Sample/ack
      -- 
    -- logger for CP element group d_block_daemon_CP_3326_elements(62)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and d_block_daemon_CP_3326_elements(62)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:d_block_daemon_CP_3326_elements(62) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:WPIPE_out_buf_10037_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_3594_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_out_buf_10037_inst_ack_0, ack => d_block_daemon_CP_3326_elements(62)); -- 
    -- CP-element group 63:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	61 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	8 
    -- CP-element group 63: marked-successors 
    -- CP-element group 63: 	61 
    -- CP-element group 63:  members (4) 
      -- CP-element group 63: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/$exit
      -- CP-element group 63: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/WPIPE_out_buf_10037_update_completed_
      -- CP-element group 63: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/WPIPE_out_buf_10037_Update/$exit
      -- CP-element group 63: 	 branch_block_stmt_9973/do_while_stmt_9974/do_while_stmt_9974_loop_body/WPIPE_out_buf_10037_Update/ack
      -- 
    -- logger for CP element group d_block_daemon_CP_3326_elements(63)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and d_block_daemon_CP_3326_elements(63)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:d_block_daemon_CP_3326_elements(63) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:WPIPE_out_buf_10037_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_3599_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_out_buf_10037_inst_ack_1, ack => d_block_daemon_CP_3326_elements(63)); -- 
    -- CP-element group 64:  transition  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	7 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	65 
    -- CP-element group 64:  members (1) 
      -- CP-element group 64: 	 branch_block_stmt_9973/do_while_stmt_9974/loop_exit/$entry
      -- 
    -- logger for CP element group d_block_daemon_CP_3326_elements(64)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and d_block_daemon_CP_3326_elements(64)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:d_block_daemon_CP_3326_elements(64) fired."); 
        -- 
      end if; --
    end process; 
    d_block_daemon_CP_3326_elements(64) <= d_block_daemon_CP_3326_elements(7);
    -- CP-element group 65:  transition  input  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	64 
    -- CP-element group 65: successors 
    -- CP-element group 65:  members (2) 
      -- CP-element group 65: 	 branch_block_stmt_9973/do_while_stmt_9974/loop_exit/$exit
      -- CP-element group 65: 	 branch_block_stmt_9973/do_while_stmt_9974/loop_exit/ack
      -- 
    -- logger for CP element group d_block_daemon_CP_3326_elements(65)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and d_block_daemon_CP_3326_elements(65)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:d_block_daemon_CP_3326_elements(65) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:do_while_stmt_9974_branch_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_3603_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_9974_branch_ack_0, ack => d_block_daemon_CP_3326_elements(65)); -- 
    -- CP-element group 66:  transition  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	7 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66:  members (1) 
      -- CP-element group 66: 	 branch_block_stmt_9973/do_while_stmt_9974/loop_taken/$entry
      -- 
    -- logger for CP element group d_block_daemon_CP_3326_elements(66)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and d_block_daemon_CP_3326_elements(66)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:d_block_daemon_CP_3326_elements(66) fired."); 
        -- 
      end if; --
    end process; 
    d_block_daemon_CP_3326_elements(66) <= d_block_daemon_CP_3326_elements(7);
    -- CP-element group 67:  transition  input  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67:  members (2) 
      -- CP-element group 67: 	 branch_block_stmt_9973/do_while_stmt_9974/loop_taken/$exit
      -- CP-element group 67: 	 branch_block_stmt_9973/do_while_stmt_9974/loop_taken/ack
      -- 
    -- logger for CP element group d_block_daemon_CP_3326_elements(67)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and d_block_daemon_CP_3326_elements(67)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:d_block_daemon_CP_3326_elements(67) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:do_while_stmt_9974_branch_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_3607_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_9974_branch_ack_1, ack => d_block_daemon_CP_3326_elements(67)); -- 
    -- CP-element group 68:  transition  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	5 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	2 
    -- CP-element group 68:  members (1) 
      -- CP-element group 68: 	 branch_block_stmt_9973/do_while_stmt_9974/$exit
      -- 
    -- logger for CP element group d_block_daemon_CP_3326_elements(68)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and d_block_daemon_CP_3326_elements(68)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:d_block_daemon_CP_3326_elements(68) fired."); 
        -- 
      end if; --
    end process; 
    d_block_daemon_CP_3326_elements(68) <= d_block_daemon_CP_3326_elements(5);
    -- CP-element group 69:  transition  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	2 
    -- CP-element group 69: successors 
    -- CP-element group 69:  members (2) 
      -- CP-element group 69: 	 $exit
      -- CP-element group 69: 	 branch_block_stmt_9973/$exit
      -- 
    -- logger for CP element group d_block_daemon_CP_3326_elements(69)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and d_block_daemon_CP_3326_elements(69)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:d_block_daemon:CP:d_block_daemon_CP_3326_elements(69) fired."); 
        -- 
      end if; --
    end process; 
    d_block_daemon_CP_3326_elements(69) <= d_block_daemon_CP_3326_elements(2);
    do_while_stmt_9974_terminator_3608: loop_terminator -- 
      generic map (max_iterations_in_flight =>10) 
      port map(loop_body_exit => d_block_daemon_CP_3326_elements(8),loop_continue => d_block_daemon_CP_3326_elements(67),loop_terminate => d_block_daemon_CP_3326_elements(65),loop_back => d_block_daemon_CP_3326_elements(6),loop_exit => d_block_daemon_CP_3326_elements(5),clk => clk, reset => reset); -- 
    entry_tmerge_3351_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= d_block_daemon_CP_3326_elements(9);
        preds(1)  <= d_block_daemon_CP_3326_elements(10);
        entry_tmerge_3351 : transition_merge -- 
          port map (preds => preds, symbol_out => d_block_daemon_CP_3326_elements(11));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_K0_10033_wire_constant : std_logic_vector(127 downto 0);
    signal R_K10_9981_wire_constant : std_logic_vector(127 downto 0);
    signal R_K1_10028_wire_constant : std_logic_vector(127 downto 0);
    signal R_K2_10023_wire_constant : std_logic_vector(127 downto 0);
    signal R_K3_10018_wire_constant : std_logic_vector(127 downto 0);
    signal R_K4_10013_wire_constant : std_logic_vector(127 downto 0);
    signal R_K5_10008_wire_constant : std_logic_vector(127 downto 0);
    signal R_K6_10003_wire_constant : std_logic_vector(127 downto 0);
    signal R_K7_9998_wire_constant : std_logic_vector(127 downto 0);
    signal R_K8_9993_wire_constant : std_logic_vector(127 downto 0);
    signal R_K9_9988_wire_constant : std_logic_vector(127 downto 0);
    signal R_LAST_9989_wire_constant : std_logic_vector(0 downto 0);
    signal R_NOT_LAST_10004_wire_constant : std_logic_vector(0 downto 0);
    signal R_NOT_LAST_10009_wire_constant : std_logic_vector(0 downto 0);
    signal R_NOT_LAST_10014_wire_constant : std_logic_vector(0 downto 0);
    signal R_NOT_LAST_10019_wire_constant : std_logic_vector(0 downto 0);
    signal R_NOT_LAST_10024_wire_constant : std_logic_vector(0 downto 0);
    signal R_NOT_LAST_10029_wire_constant : std_logic_vector(0 downto 0);
    signal R_NOT_LAST_10034_wire_constant : std_logic_vector(0 downto 0);
    signal R_NOT_LAST_9994_wire_constant : std_logic_vector(0 downto 0);
    signal R_NOT_LAST_9999_wire_constant : std_logic_vector(0 downto 0);
    signal in128_9978 : std_logic_vector(127 downto 0);
    signal konst_10041_wire_constant : std_logic_vector(0 downto 0);
    signal round_S0_10036 : std_logic_vector(127 downto 0);
    signal round_S10_9983 : std_logic_vector(127 downto 0);
    signal round_S10_9984_delayed_1_9986 : std_logic_vector(127 downto 0);
    signal round_S1_10031 : std_logic_vector(127 downto 0);
    signal round_S2_10026 : std_logic_vector(127 downto 0);
    signal round_S3_10021 : std_logic_vector(127 downto 0);
    signal round_S4_10016 : std_logic_vector(127 downto 0);
    signal round_S5_10011 : std_logic_vector(127 downto 0);
    signal round_S6_10006 : std_logic_vector(127 downto 0);
    signal round_S7_10001 : std_logic_vector(127 downto 0);
    signal round_S8_9996 : std_logic_vector(127 downto 0);
    signal round_S9_9991 : std_logic_vector(127 downto 0);
    signal xxd_block_daemonxxK0 : std_logic_vector(127 downto 0);
    signal xxd_block_daemonxxK1 : std_logic_vector(127 downto 0);
    signal xxd_block_daemonxxK10 : std_logic_vector(127 downto 0);
    signal xxd_block_daemonxxK2 : std_logic_vector(127 downto 0);
    signal xxd_block_daemonxxK3 : std_logic_vector(127 downto 0);
    signal xxd_block_daemonxxK4 : std_logic_vector(127 downto 0);
    signal xxd_block_daemonxxK5 : std_logic_vector(127 downto 0);
    signal xxd_block_daemonxxK6 : std_logic_vector(127 downto 0);
    signal xxd_block_daemonxxK7 : std_logic_vector(127 downto 0);
    signal xxd_block_daemonxxK8 : std_logic_vector(127 downto 0);
    signal xxd_block_daemonxxK9 : std_logic_vector(127 downto 0);
    signal xxd_block_daemonxxLAST : std_logic_vector(0 downto 0);
    signal xxd_block_daemonxxNOT_LAST : std_logic_vector(0 downto 0);
    signal xxd_block_daemonxxRConstant_1 : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    R_K0_10033_wire_constant <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    R_K10_9981_wire_constant <= "10110100111011110101101111001011001111101001001011100010000100010010001111101001010100011100111101101111100011110001100010001110";
    R_K1_10028_wire_constant <= "01100010011000110110001101100011011000100110001101100011011000110110001001100011011000110110001101100010011000110110001101100011";
    R_K2_10023_wire_constant <= "10011011100110001001100011001001111110011111101111111011101010101001101110011000100110001100100111111001111110111111101110101010";
    R_K3_10018_wire_constant <= "10010000100101110011010001010000011010010110110011001111111110101111001011110100010101110011001100001011000011111010110010011001";
    R_K4_10013_wire_constant <= "11101110000001101101101001111011100001110110101000010101100000010111010110011110010000101011001001111110100100011110111000101011";
    R_K5_10008_wire_constant <= "01111111001011100010101110001000111110000100010000111110000010011000110111011010011111001011101111110011010010111001001010010000";
    R_K6_10003_wire_constant <= "11101100011000010100101110000101000101000010010101110101100011001001100111111111000010010011011101101010101101001001101110100111";
    R_K7_9998_wire_constant <= "00100001011101010001011110000111001101010101000001100010000010111010110010101111011010110011110011000110000110111111000010011011";
    R_K8_9993_wire_constant <= "00001110111110010000001100110011001110111010100101100001001110001001011100000110000010100000010001010001000111011111101010011111";
    R_K9_9988_wire_constant <= "10110001110101001101100011100010100010100111110110111001110110100001110101111011101100111101111001001100011001100100100101000001";
    R_LAST_9989_wire_constant <= "1";
    R_NOT_LAST_10004_wire_constant <= "0";
    R_NOT_LAST_10009_wire_constant <= "0";
    R_NOT_LAST_10014_wire_constant <= "0";
    R_NOT_LAST_10019_wire_constant <= "0";
    R_NOT_LAST_10024_wire_constant <= "0";
    R_NOT_LAST_10029_wire_constant <= "0";
    R_NOT_LAST_10034_wire_constant <= "0";
    R_NOT_LAST_9994_wire_constant <= "0";
    R_NOT_LAST_9999_wire_constant <= "0";
    konst_10041_wire_constant <= "1";
    xxd_block_daemonxxK0 <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    xxd_block_daemonxxK1 <= "01100010011000110110001101100011011000100110001101100011011000110110001001100011011000110110001101100010011000110110001101100011";
    xxd_block_daemonxxK10 <= "10110100111011110101101111001011001111101001001011100010000100010010001111101001010100011100111101101111100011110001100010001110";
    xxd_block_daemonxxK2 <= "10011011100110001001100011001001111110011111101111111011101010101001101110011000100110001100100111111001111110111111101110101010";
    xxd_block_daemonxxK3 <= "10010000100101110011010001010000011010010110110011001111111110101111001011110100010101110011001100001011000011111010110010011001";
    xxd_block_daemonxxK4 <= "11101110000001101101101001111011100001110110101000010101100000010111010110011110010000101011001001111110100100011110111000101011";
    xxd_block_daemonxxK5 <= "01111111001011100010101110001000111110000100010000111110000010011000110111011010011111001011101111110011010010111001001010010000";
    xxd_block_daemonxxK6 <= "11101100011000010100101110000101000101000010010101110101100011001001100111111111000010010011011101101010101101001001101110100111";
    xxd_block_daemonxxK7 <= "00100001011101010001011110000111001101010101000001100010000010111010110010101111011010110011110011000110000110111111000010011011";
    xxd_block_daemonxxK8 <= "00001110111110010000001100110011001110111010100101100001001110001001011100000110000010100000010001010001000111011111101010011111";
    xxd_block_daemonxxK9 <= "10110001110101001101100011100010100010100111110110111001110110100001110101111011101100111101111001001100011001100100100101000001";
    xxd_block_daemonxxLAST <= "1";
    xxd_block_daemonxxNOT_LAST <= "0";
    xxd_block_daemonxxRConstant_1 <= "00000001";
    -- logger for split-operator W_round_S10_9984_delayed_1_9984_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if W_round_S10_9984_delayed_1_9984_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:d_block_daemon:DP:W_round_S10_9984_delayed_1_9984_inst:started:   inputs: " & " round_S10_9983 = "& Convert_SLV_To_Hex_String(round_S10_9983));
          --
        end if; 
        if W_round_S10_9984_delayed_1_9984_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:d_block_daemon:DP:W_round_S10_9984_delayed_1_9984_inst:finished:  outputs: " & " round_S10_9984_delayed_1_9986= "  & Convert_SLV_To_Hex_String(round_S10_9984_delayed_1_9986));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    W_round_S10_9984_delayed_1_9984_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_round_S10_9984_delayed_1_9984_inst_req_0;
      W_round_S10_9984_delayed_1_9984_inst_ack_0<= wack(0);
      rreq(0) <= W_round_S10_9984_delayed_1_9984_inst_req_1;
      W_round_S10_9984_delayed_1_9984_inst_ack_1<= rack(0);
      W_round_S10_9984_delayed_1_9984_inst : InterlockBuffer generic map ( -- 
        name => "W_round_S10_9984_delayed_1_9984_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 128,
        out_data_width => 128,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => round_S10_9983,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => round_S10_9984_delayed_1_9986,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_9974_branch_req_0," req0 do_while_stmt_9974_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_9974_branch_ack_0," ack0 do_while_stmt_9974_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_9974_branch_ack_1," ack1 do_while_stmt_9974_branch");
    do_while_stmt_9974_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= konst_10041_wire_constant;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_9974_branch_req_0,
          ack0 => do_while_stmt_9974_branch_ack_0,
          ack1 => do_while_stmt_9974_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- logger for split-operator XOR_u128_u128_9982_inst flow-through 
    process(round_S10_9983) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:d_block_daemon:DP:XOR_u128_u128_9982_inst:flowthrough inputs: " & " in128_9978 = "& Convert_SLV_To_Hex_String(in128_9978) & " R_K10_9981_wire_constant = "& Convert_SLV_To_Hex_String(R_K10_9981_wire_constant) & " outputs:" & " round_S10_9983= "  & Convert_SLV_To_Hex_String(round_S10_9983));
      --
    end process; 
    -- binary operator XOR_u128_u128_9982_inst
    process(in128_9978) -- 
      variable tmp_var : std_logic_vector(127 downto 0); -- 
    begin -- 
      ApIntXor_proc(in128_9978, R_K10_9981_wire_constant, tmp_var);
      round_S10_9983 <= tmp_var; -- 
    end process;
    -- logger for split-operator RPIPE_in_buf_9977_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if RPIPE_in_buf_9977_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:d_block_daemon:DP:RPIPE_in_buf_9977_inst:started:   PipeRead from in_buf inputs: " & " no-guard, no-inputs ");
          --
        end if; 
        if RPIPE_in_buf_9977_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:d_block_daemon:DP:RPIPE_in_buf_9977_inst:finished:  outputs: " & " in128_9978= "  & Convert_SLV_To_Hex_String(in128_9978));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared inport operator group (0) : RPIPE_in_buf_9977_inst 
    InportGroup0: Block -- 
      signal data_out: std_logic_vector(127 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_in_buf_9977_inst_req_0;
      RPIPE_in_buf_9977_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_in_buf_9977_inst_req_1;
      RPIPE_in_buf_9977_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      in128_9978 <= data_out(127 downto 0);
      in_buf_read_0: InputPortRevised -- 
        generic map ( name => "in_buf_read_0", data_width => 128,  num_reqs => 1,  output_buffering => outBUFs,   no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => in_buf_pipe_read_req(0),
          oack => in_buf_pipe_read_ack(0),
          odata => in_buf_pipe_read_data(127 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- logger for split-operator WPIPE_out_buf_10037_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if WPIPE_out_buf_10037_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:d_block_daemon:DP:WPIPE_out_buf_10037_inst:started:   PipeWrite to out_buf inputs: " & " round_S0_10036 = "& Convert_SLV_To_Hex_String(round_S0_10036));
          --
        end if; 
        if WPIPE_out_buf_10037_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:d_block_daemon:DP:WPIPE_out_buf_10037_inst:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared outport operator group (0) : WPIPE_out_buf_10037_inst 
    OutportGroup0: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_out_buf_10037_inst_req_0;
      WPIPE_out_buf_10037_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_out_buf_10037_inst_req_1;
      WPIPE_out_buf_10037_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      data_in <= round_S0_10036;
      out_buf_write_0: OutputPortRevised -- 
        generic map ( name => "out_buf", data_width => 128, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => out_buf_pipe_write_req(0),
          oack => out_buf_pipe_write_ack(0),
          odata => out_buf_pipe_write_data(127 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- logger for split-operator call_stmt_10001_call
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if call_stmt_10001_call_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:d_block_daemon:DP:call_stmt_10001_call:started:  Call to module dec_round inputs: " & " round_S8_9996 = "& Convert_SLV_To_Hex_String(round_S8_9996) & " R_K7_9998_wire_constant = "& Convert_SLV_To_Hex_String(R_K7_9998_wire_constant) & " R_NOT_LAST_9999_wire_constant = "& Convert_SLV_To_Hex_String(R_NOT_LAST_9999_wire_constant));
          --
        end if; 
        if call_stmt_10001_call_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:d_block_daemon:DP:call_stmt_10001_call:finished:  outputs: " & " round_S7_10001= "  & Convert_SLV_To_Hex_String(round_S7_10001));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    call_stmt_10001_call_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= call_stmt_10001_call_req_0;
      call_stmt_10001_call_ack_0<= sample_ack(0);
      update_req(0) <= call_stmt_10001_call_req_1;
      call_stmt_10001_call_ack_1<= update_ack(0);
      call_stmt_10001_call: dec_round_Operator  port map ( -- 
        sample_req => sample_req(0), 
        sample_ack => sample_ack(0), 
        update_req => update_req(0), 
        update_ack => update_ack(0), 
        round_in => round_S8_9996,
        key_in => R_K7_9998_wire_constant,
        l_round => R_NOT_LAST_9999_wire_constant,
        round_out => round_S7_10001,
        clk => clk, reset => reset  
        -- 
      );-- 
    end block;
    -- logger for split-operator call_stmt_10006_call
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if call_stmt_10006_call_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:d_block_daemon:DP:call_stmt_10006_call:started:  Call to module dec_round inputs: " & " round_S7_10001 = "& Convert_SLV_To_Hex_String(round_S7_10001) & " R_K6_10003_wire_constant = "& Convert_SLV_To_Hex_String(R_K6_10003_wire_constant) & " R_NOT_LAST_10004_wire_constant = "& Convert_SLV_To_Hex_String(R_NOT_LAST_10004_wire_constant));
          --
        end if; 
        if call_stmt_10006_call_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:d_block_daemon:DP:call_stmt_10006_call:finished:  outputs: " & " round_S6_10006= "  & Convert_SLV_To_Hex_String(round_S6_10006));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    call_stmt_10006_call_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= call_stmt_10006_call_req_0;
      call_stmt_10006_call_ack_0<= sample_ack(0);
      update_req(0) <= call_stmt_10006_call_req_1;
      call_stmt_10006_call_ack_1<= update_ack(0);
      call_stmt_10006_call: dec_round_Operator  port map ( -- 
        sample_req => sample_req(0), 
        sample_ack => sample_ack(0), 
        update_req => update_req(0), 
        update_ack => update_ack(0), 
        round_in => round_S7_10001,
        key_in => R_K6_10003_wire_constant,
        l_round => R_NOT_LAST_10004_wire_constant,
        round_out => round_S6_10006,
        clk => clk, reset => reset  
        -- 
      );-- 
    end block;
    -- logger for split-operator call_stmt_10011_call
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if call_stmt_10011_call_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:d_block_daemon:DP:call_stmt_10011_call:started:  Call to module dec_round inputs: " & " round_S6_10006 = "& Convert_SLV_To_Hex_String(round_S6_10006) & " R_K5_10008_wire_constant = "& Convert_SLV_To_Hex_String(R_K5_10008_wire_constant) & " R_NOT_LAST_10009_wire_constant = "& Convert_SLV_To_Hex_String(R_NOT_LAST_10009_wire_constant));
          --
        end if; 
        if call_stmt_10011_call_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:d_block_daemon:DP:call_stmt_10011_call:finished:  outputs: " & " round_S5_10011= "  & Convert_SLV_To_Hex_String(round_S5_10011));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    call_stmt_10011_call_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= call_stmt_10011_call_req_0;
      call_stmt_10011_call_ack_0<= sample_ack(0);
      update_req(0) <= call_stmt_10011_call_req_1;
      call_stmt_10011_call_ack_1<= update_ack(0);
      call_stmt_10011_call: dec_round_Operator  port map ( -- 
        sample_req => sample_req(0), 
        sample_ack => sample_ack(0), 
        update_req => update_req(0), 
        update_ack => update_ack(0), 
        round_in => round_S6_10006,
        key_in => R_K5_10008_wire_constant,
        l_round => R_NOT_LAST_10009_wire_constant,
        round_out => round_S5_10011,
        clk => clk, reset => reset  
        -- 
      );-- 
    end block;
    -- logger for split-operator call_stmt_10016_call
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if call_stmt_10016_call_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:d_block_daemon:DP:call_stmt_10016_call:started:  Call to module dec_round inputs: " & " round_S5_10011 = "& Convert_SLV_To_Hex_String(round_S5_10011) & " R_K4_10013_wire_constant = "& Convert_SLV_To_Hex_String(R_K4_10013_wire_constant) & " R_NOT_LAST_10014_wire_constant = "& Convert_SLV_To_Hex_String(R_NOT_LAST_10014_wire_constant));
          --
        end if; 
        if call_stmt_10016_call_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:d_block_daemon:DP:call_stmt_10016_call:finished:  outputs: " & " round_S4_10016= "  & Convert_SLV_To_Hex_String(round_S4_10016));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    call_stmt_10016_call_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= call_stmt_10016_call_req_0;
      call_stmt_10016_call_ack_0<= sample_ack(0);
      update_req(0) <= call_stmt_10016_call_req_1;
      call_stmt_10016_call_ack_1<= update_ack(0);
      call_stmt_10016_call: dec_round_Operator  port map ( -- 
        sample_req => sample_req(0), 
        sample_ack => sample_ack(0), 
        update_req => update_req(0), 
        update_ack => update_ack(0), 
        round_in => round_S5_10011,
        key_in => R_K4_10013_wire_constant,
        l_round => R_NOT_LAST_10014_wire_constant,
        round_out => round_S4_10016,
        clk => clk, reset => reset  
        -- 
      );-- 
    end block;
    -- logger for split-operator call_stmt_10021_call
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if call_stmt_10021_call_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:d_block_daemon:DP:call_stmt_10021_call:started:  Call to module dec_round inputs: " & " round_S4_10016 = "& Convert_SLV_To_Hex_String(round_S4_10016) & " R_K3_10018_wire_constant = "& Convert_SLV_To_Hex_String(R_K3_10018_wire_constant) & " R_NOT_LAST_10019_wire_constant = "& Convert_SLV_To_Hex_String(R_NOT_LAST_10019_wire_constant));
          --
        end if; 
        if call_stmt_10021_call_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:d_block_daemon:DP:call_stmt_10021_call:finished:  outputs: " & " round_S3_10021= "  & Convert_SLV_To_Hex_String(round_S3_10021));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    call_stmt_10021_call_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= call_stmt_10021_call_req_0;
      call_stmt_10021_call_ack_0<= sample_ack(0);
      update_req(0) <= call_stmt_10021_call_req_1;
      call_stmt_10021_call_ack_1<= update_ack(0);
      call_stmt_10021_call: dec_round_Operator  port map ( -- 
        sample_req => sample_req(0), 
        sample_ack => sample_ack(0), 
        update_req => update_req(0), 
        update_ack => update_ack(0), 
        round_in => round_S4_10016,
        key_in => R_K3_10018_wire_constant,
        l_round => R_NOT_LAST_10019_wire_constant,
        round_out => round_S3_10021,
        clk => clk, reset => reset  
        -- 
      );-- 
    end block;
    -- logger for split-operator call_stmt_10026_call
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if call_stmt_10026_call_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:d_block_daemon:DP:call_stmt_10026_call:started:  Call to module dec_round inputs: " & " round_S3_10021 = "& Convert_SLV_To_Hex_String(round_S3_10021) & " R_K2_10023_wire_constant = "& Convert_SLV_To_Hex_String(R_K2_10023_wire_constant) & " R_NOT_LAST_10024_wire_constant = "& Convert_SLV_To_Hex_String(R_NOT_LAST_10024_wire_constant));
          --
        end if; 
        if call_stmt_10026_call_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:d_block_daemon:DP:call_stmt_10026_call:finished:  outputs: " & " round_S2_10026= "  & Convert_SLV_To_Hex_String(round_S2_10026));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    call_stmt_10026_call_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= call_stmt_10026_call_req_0;
      call_stmt_10026_call_ack_0<= sample_ack(0);
      update_req(0) <= call_stmt_10026_call_req_1;
      call_stmt_10026_call_ack_1<= update_ack(0);
      call_stmt_10026_call: dec_round_Operator  port map ( -- 
        sample_req => sample_req(0), 
        sample_ack => sample_ack(0), 
        update_req => update_req(0), 
        update_ack => update_ack(0), 
        round_in => round_S3_10021,
        key_in => R_K2_10023_wire_constant,
        l_round => R_NOT_LAST_10024_wire_constant,
        round_out => round_S2_10026,
        clk => clk, reset => reset  
        -- 
      );-- 
    end block;
    -- logger for split-operator call_stmt_10031_call
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if call_stmt_10031_call_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:d_block_daemon:DP:call_stmt_10031_call:started:  Call to module dec_round inputs: " & " round_S2_10026 = "& Convert_SLV_To_Hex_String(round_S2_10026) & " R_K1_10028_wire_constant = "& Convert_SLV_To_Hex_String(R_K1_10028_wire_constant) & " R_NOT_LAST_10029_wire_constant = "& Convert_SLV_To_Hex_String(R_NOT_LAST_10029_wire_constant));
          --
        end if; 
        if call_stmt_10031_call_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:d_block_daemon:DP:call_stmt_10031_call:finished:  outputs: " & " round_S1_10031= "  & Convert_SLV_To_Hex_String(round_S1_10031));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    call_stmt_10031_call_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= call_stmt_10031_call_req_0;
      call_stmt_10031_call_ack_0<= sample_ack(0);
      update_req(0) <= call_stmt_10031_call_req_1;
      call_stmt_10031_call_ack_1<= update_ack(0);
      call_stmt_10031_call: dec_round_Operator  port map ( -- 
        sample_req => sample_req(0), 
        sample_ack => sample_ack(0), 
        update_req => update_req(0), 
        update_ack => update_ack(0), 
        round_in => round_S2_10026,
        key_in => R_K1_10028_wire_constant,
        l_round => R_NOT_LAST_10029_wire_constant,
        round_out => round_S1_10031,
        clk => clk, reset => reset  
        -- 
      );-- 
    end block;
    -- logger for split-operator call_stmt_10036_call
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if call_stmt_10036_call_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:d_block_daemon:DP:call_stmt_10036_call:started:  Call to module dec_round inputs: " & " round_S1_10031 = "& Convert_SLV_To_Hex_String(round_S1_10031) & " R_K0_10033_wire_constant = "& Convert_SLV_To_Hex_String(R_K0_10033_wire_constant) & " R_NOT_LAST_10034_wire_constant = "& Convert_SLV_To_Hex_String(R_NOT_LAST_10034_wire_constant));
          --
        end if; 
        if call_stmt_10036_call_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:d_block_daemon:DP:call_stmt_10036_call:finished:  outputs: " & " round_S0_10036= "  & Convert_SLV_To_Hex_String(round_S0_10036));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    call_stmt_10036_call_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= call_stmt_10036_call_req_0;
      call_stmt_10036_call_ack_0<= sample_ack(0);
      update_req(0) <= call_stmt_10036_call_req_1;
      call_stmt_10036_call_ack_1<= update_ack(0);
      call_stmt_10036_call: dec_round_Operator  port map ( -- 
        sample_req => sample_req(0), 
        sample_ack => sample_ack(0), 
        update_req => update_req(0), 
        update_ack => update_ack(0), 
        round_in => round_S1_10031,
        key_in => R_K0_10033_wire_constant,
        l_round => R_NOT_LAST_10034_wire_constant,
        round_out => round_S0_10036,
        clk => clk, reset => reset  
        -- 
      );-- 
    end block;
    -- logger for split-operator call_stmt_9991_call
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if call_stmt_9991_call_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:d_block_daemon:DP:call_stmt_9991_call:started:  Call to module dec_round inputs: " & " round_S10_9984_delayed_1_9986 = "& Convert_SLV_To_Hex_String(round_S10_9984_delayed_1_9986) & " R_K9_9988_wire_constant = "& Convert_SLV_To_Hex_String(R_K9_9988_wire_constant) & " R_LAST_9989_wire_constant = "& Convert_SLV_To_Hex_String(R_LAST_9989_wire_constant));
          --
        end if; 
        if call_stmt_9991_call_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:d_block_daemon:DP:call_stmt_9991_call:finished:  outputs: " & " round_S9_9991= "  & Convert_SLV_To_Hex_String(round_S9_9991));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    call_stmt_9991_call_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= call_stmt_9991_call_req_0;
      call_stmt_9991_call_ack_0<= sample_ack(0);
      update_req(0) <= call_stmt_9991_call_req_1;
      call_stmt_9991_call_ack_1<= update_ack(0);
      call_stmt_9991_call: dec_round_Operator  port map ( -- 
        sample_req => sample_req(0), 
        sample_ack => sample_ack(0), 
        update_req => update_req(0), 
        update_ack => update_ack(0), 
        round_in => round_S10_9984_delayed_1_9986,
        key_in => R_K9_9988_wire_constant,
        l_round => R_LAST_9989_wire_constant,
        round_out => round_S9_9991,
        clk => clk, reset => reset  
        -- 
      );-- 
    end block;
    -- logger for split-operator call_stmt_9996_call
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if call_stmt_9996_call_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:d_block_daemon:DP:call_stmt_9996_call:started:  Call to module dec_round inputs: " & " round_S9_9991 = "& Convert_SLV_To_Hex_String(round_S9_9991) & " R_K8_9993_wire_constant = "& Convert_SLV_To_Hex_String(R_K8_9993_wire_constant) & " R_NOT_LAST_9994_wire_constant = "& Convert_SLV_To_Hex_String(R_NOT_LAST_9994_wire_constant));
          --
        end if; 
        if call_stmt_9996_call_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:d_block_daemon:DP:call_stmt_9996_call:finished:  outputs: " & " round_S8_9996= "  & Convert_SLV_To_Hex_String(round_S8_9996));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    call_stmt_9996_call_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= call_stmt_9996_call_req_0;
      call_stmt_9996_call_ack_0<= sample_ack(0);
      update_req(0) <= call_stmt_9996_call_req_1;
      call_stmt_9996_call_ack_1<= update_ack(0);
      call_stmt_9996_call: dec_round_Operator  port map ( -- 
        sample_req => sample_req(0), 
        sample_ack => sample_ack(0), 
        update_req => update_req(0), 
        update_ack => update_ack(0), 
        round_in => round_S9_9991,
        key_in => R_K8_9993_wire_constant,
        l_round => R_NOT_LAST_9994_wire_constant,
        round_out => round_S8_9996,
        clk => clk, reset => reset  
        -- 
      );-- 
    end block;
    -- 
  end Block; -- data_path
  -- 
end d_block_daemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library GhdlLink;
use GhdlLink.LogUtilities.all;
library work;
use work.ahir_system_global_package.all;
entity dec_round_Operator is -- 
  port ( -- 
    sample_req: in boolean;
    sample_ack: out boolean;
    update_req: in boolean;
    update_ack: out boolean;
    round_in : in  std_logic_vector(127 downto 0);
    key_in : in  std_logic_vector(127 downto 0);
    l_round : in  std_logic_vector(0 downto 0);
    round_out : out  std_logic_vector(127 downto 0);
    clk, reset: in std_logic
    -- 
  );
  -- 
end entity dec_round_Operator;
architecture dec_round_Operator_arch of dec_round_Operator is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal update_ack_symbol: Boolean;
  signal default_zero_sig: std_logic;
  -- input port buffer signals
  signal round_in_buffer :  std_logic_vector(127 downto 0);
  signal round_in_update_enable: Boolean;
  signal round_in_update_enable_unmarked: Boolean;
  signal key_in_buffer :  std_logic_vector(127 downto 0);
  signal key_in_update_enable: Boolean;
  signal key_in_update_enable_unmarked: Boolean;
  signal l_round_buffer :  std_logic_vector(0 downto 0);
  signal l_round_update_enable: Boolean;
  signal l_round_update_enable_unmarked: Boolean;
  -- output port buffer signals
  signal round_out_buffer :  std_logic_vector(127 downto 0);
  signal round_out_update_enable: Boolean;
  signal dec_round_CP_192_start: Boolean;
  signal dec_round_CP_192_symbol: Boolean;
  signal cp_all_inputs_sampled: Boolean;
  -- volatile/operator module components. 
  component Inv_Sbox_2_Volatile is -- 
    port ( -- 
      clk, reset: in std_logic; 
      s_in : in  std_logic_vector(7 downto 0);
      s_out : out  std_logic_vector(7 downto 0)-- 
    );
    -- 
  end component; 
  component Inv_Sbox_1_Volatile is -- 
    port ( -- 
      clk, reset: in std_logic; 
      s_in : in  std_logic_vector(7 downto 0);
      s_out : out  std_logic_vector(7 downto 0)-- 
    );
    -- 
  end component; 
  component Inv_Sbox_3_Volatile is -- 
    port ( -- 
      clk, reset: in std_logic; 
      s_in : in  std_logic_vector(7 downto 0);
      s_out : out  std_logic_vector(7 downto 0)-- 
    );
    -- 
  end component; 
  component Inv_Sbox_4_Volatile is -- 
    port ( -- 
      clk, reset: in std_logic; 
      s_in : in  std_logic_vector(7 downto 0);
      s_out : out  std_logic_vector(7 downto 0)-- 
    );
    -- 
  end component; 
  component MUL2_Volatile is -- 
    port ( -- 
      clk, reset: in std_logic; 
      mul_in : in  std_logic_vector(7 downto 0);
      mul_out : out  std_logic_vector(7 downto 0)-- 
    );
    -- 
  end component; 
  -- links between control-path and data-path
  signal XOR_u128_u128_9927_inst_ack_1 : boolean;
  signal XOR_u128_u128_9927_inst_req_1 : boolean;
  signal XOR_u128_u128_9927_inst_ack_0 : boolean;
  signal XOR_u128_u128_9927_inst_req_0 : boolean;
  signal global_clock_cycle_count: integer := 0;
  -- 
begin --  
  ---------------------------------------------------------- 
  process(clk)  
  begin -- 
    if(clk'event and clk = '1') then -- 
      if(reset = '1') then -- 
        global_clock_cycle_count <= 0; --
      else -- 
        global_clock_cycle_count <= global_clock_cycle_count + 1; -- 
      end if; --
    end if; --
  end process;
  ---------------------------------------------------------- 
  sample_ack <= dec_round_CP_192_symbol;
  -- input handling ------------------------------------------------
  round_in_buffer <= round_in;
  key_in_buffer <= key_in;
  l_round_buffer <= l_round;
  dec_round_CP_192_start <= sample_req;
  -- output handling  -------------------------------------------------------
  round_out <= round_out_buffer;
  round_out_update_enable <= update_req;
  update_ack_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 22) := "update_ack_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= dec_round_CP_192_symbol & update_req;
    gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => update_ack_symbol, clk => clk, reset => reset); --
  end block;
  -- update ack. 
  update_ack <= update_ack_symbol;
  --- logging ------------------------------------------------------
  LogCPEvent(clk,reset,global_clock_cycle_count,dec_round_CP_192_start,"dec_round cp_entry_symbol ");
  LogCPEvent(clk,reset,global_clock_cycle_count,dec_round_CP_192_symbol, "dec_round cp_exit_symbol ");
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  dec_round_CP_192: Block -- control-path 
    signal dec_round_CP_192_elements: BooleanArray(2 downto 0);
    -- 
  begin -- 
    dec_round_CP_192_elements(0) <= dec_round_CP_192_start;
    dec_round_CP_192_symbol <= dec_round_CP_192_elements(2);
    -- CP-element group 0:  join  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (2852) 
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9329_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9353_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISd_9340_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9321_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9353_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISd_9340_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9329_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9349_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9333_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9325_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS02_9357_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9337_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISd_9340_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9341_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS06_9369_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9321_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9333_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISc_9320_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9374_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9341_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISc_9324_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISc_9332_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISd_9344_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9325_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9325_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9349_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9329_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9365_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9333_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9333_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS06_9369_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS03_9360_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS04_9363_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS03_9360_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9368_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISc_9332_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS08_9375_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9337_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9345_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9345_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9337_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS02_9357_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS06_9369_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9341_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9325_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISd_9340_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9341_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS09_9378_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9345_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS00_9351_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9353_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9333_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9325_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9389_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISc_9320_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9365_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISd_9344_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9353_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS08_9375_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9345_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS10_9381_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9325_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9333_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9333_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISc_9320_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9341_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9377_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9480_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9333_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9337_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9380_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS04_9363_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS00_9351_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9325_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS05_9366_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9380_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9483_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9337_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS09_9378_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Y00_9475_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9337_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9341_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISd_9344_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9386_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISd_9344_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISc_9320_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS00_9351_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9356_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9345_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9345_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9341_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9345_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9383_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9365_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISc_9332_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9365_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9386_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9383_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9325_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9371_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9345_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISc_9332_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9321_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9374_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS00_9351_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS05_9366_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS04_9363_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9329_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS01_9354_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS01_9354_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9368_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9333_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9383_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9345_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9374_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS01_9354_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9337_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9345_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS12_9387_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9329_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9368_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS10_9381_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9341_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS01_9354_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9359_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9368_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9362_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9341_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9345_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS02_9357_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9329_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9329_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9345_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9359_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9349_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9359_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9377_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS03_9360_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9386_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Y01_9478_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9374_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9333_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9349_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9389_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS11_9384_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISc_9328_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS11_9384_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9356_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISc_9328_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9359_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9349_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9377_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9341_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS03_9360_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9371_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9362_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9349_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9333_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9383_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Y00_9475_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISd_9348_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9389_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Y01_9478_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS08_9375_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9389_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9341_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISc_9328_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISd_9348_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9356_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS11_9384_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9362_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS06_9369_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9380_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS09_9378_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISd_9348_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISc_9328_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS02_9357_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISd_9348_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS07_9372_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9341_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9349_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS05_9366_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9329_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9329_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9329_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS11_9384_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9329_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS09_9378_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9333_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS10_9381_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS05_9366_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9349_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9329_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS08_9375_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9356_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9325_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9325_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9321_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9380_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9377_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS07_9372_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS07_9372_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9386_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS04_9363_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS10_9381_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Y02_9481_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS07_9372_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9371_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9371_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9498_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9337_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9530_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9498_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISd_9336_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Y13x2_9516_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISd_9336_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISc_9324_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9362_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9349_Update/cr
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9273_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9273_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9273_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9273_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_round_in_9271_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_round_in_9271_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_round_in_9271_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_round_in_9271_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISc_9324_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9321_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISd_9336_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9321_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISd_9336_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9273_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9273_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9273_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9273_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISc_9324_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9273_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9273_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9273_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9273_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9349_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9277_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9277_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9277_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9277_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_round_in_9276_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_round_in_9276_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_round_in_9276_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_round_in_9276_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9325_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9321_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9337_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9321_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9337_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9277_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9277_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9277_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9277_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9277_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9277_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9277_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9277_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9483_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9349_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9281_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9281_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9281_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9281_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_round_in_9280_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_round_in_9280_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_round_in_9280_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_round_in_9280_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9325_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9321_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9337_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9321_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9337_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9281_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9281_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9281_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9281_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9281_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9281_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9281_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9281_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9483_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9349_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9285_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9285_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9285_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9285_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_round_in_9284_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_round_in_9284_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_round_in_9284_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_round_in_9284_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9480_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9285_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9285_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9285_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9285_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9285_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9285_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9285_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9285_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Y02_9481_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9289_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9289_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9289_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9289_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISa_9288_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISa_9288_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISa_9288_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISa_9288_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Y10x2_9501_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9530_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9289_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9289_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9289_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9289_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9289_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9289_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9495_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9289_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9289_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9486_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9480_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9517_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Y13_9496_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9293_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9293_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9293_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9293_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISa_9292_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISa_9292_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISa_9292_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISa_9292_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Y01_9478_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9293_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9293_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Y12_9493_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9293_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9293_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9293_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9293_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Y12_9493_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9293_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9293_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9502_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9297_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9297_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9297_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9297_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISa_9296_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS12_9387_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9483_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISa_9296_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISa_9296_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISa_9296_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9498_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9486_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Y02_9481_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9297_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9297_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9297_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9297_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9297_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9297_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Y12_9493_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9297_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9297_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9480_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Y13_9496_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9301_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9301_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9301_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9301_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISa_9300_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISa_9300_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISa_9300_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISa_9300_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Y10x2_9501_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Y02_9481_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9486_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Y03_9484_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9301_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9301_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9301_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9301_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9301_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9301_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9301_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9301_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9305_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9305_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9305_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9305_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISb_9304_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISb_9304_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISb_9304_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISb_9304_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9305_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9305_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9305_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9305_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9305_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9305_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9305_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9305_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9309_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9309_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9309_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9309_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISb_9308_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISb_9308_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISb_9308_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISb_9308_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9309_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9309_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9309_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9309_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9309_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9309_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9309_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9309_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9313_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9313_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9313_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9313_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISb_9312_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISb_9312_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISb_9312_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISb_9312_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9313_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9313_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9313_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9313_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9313_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9313_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9313_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9313_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9317_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9317_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9317_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9317_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISb_9316_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISb_9316_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISb_9316_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISb_9316_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9317_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9317_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9317_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9317_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9317_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9317_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9317_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9317_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9321_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/slice_9321_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS12_9387_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS12_9387_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Y01_9478_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS12x2_9451_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9630_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9392_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9392_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9392_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9392_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS13_9390_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS13_9390_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS13_9390_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS13_9390_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9395_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9395_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9395_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9395_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS14_9393_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS14_9393_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS14_9393_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS14_9393_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9398_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9398_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9398_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9398_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS15_9396_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS15_9396_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS15_9396_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS15_9396_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9406_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9406_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9406_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9406_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9402_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9402_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9402_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9402_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS00_9400_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS00_9400_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS00_9400_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS00_9400_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS01_9401_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS01_9401_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS01_9401_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS01_9401_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9402_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9402_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9402_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9402_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9402_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9402_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9402_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9402_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9405_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9405_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9405_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9405_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS02_9403_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS02_9403_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS02_9403_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS02_9403_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS03_9404_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS03_9404_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS03_9404_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS03_9404_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9405_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9405_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9405_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9405_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9405_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9405_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9405_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9405_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9406_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9406_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9406_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9406_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9406_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9406_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9406_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9406_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9415_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9415_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9415_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9415_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9411_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9411_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9411_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9411_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS04_9409_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS04_9409_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS04_9409_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS04_9409_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Y01x2_9505_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Y13x2_9516_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Y13x2_9516_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS05_9410_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS05_9410_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS05_9410_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS05_9410_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Y10x2_9501_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Y01x2_9505_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Y13x2_9516_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Y03x2_9515_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Y03x2_9515_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Y03x2_9515_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9411_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9411_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9495_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9411_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9411_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9411_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9411_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9495_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9411_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9411_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Y03x2_9515_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9530_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Wc0_9533_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Wc0_9533_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Z2_9525_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Z2_9525_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9414_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9414_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9414_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9414_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS06_9412_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS06_9412_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS06_9412_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS06_9412_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Y00x2_9500_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Y01x2_9505_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9517_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9517_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS07_9413_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS07_9413_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS07_9413_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS07_9413_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Y00x2_9500_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Y01x2_9505_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9517_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9517_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9512_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9512_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9414_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9414_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9495_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9414_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9414_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9414_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9414_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Y11_9490_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9414_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9414_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9512_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Z2_9525_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Wc0_9533_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Wc0_9533_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Z2_9525_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9527_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9527_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9527_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9415_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9415_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Y11_9490_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9415_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9415_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9415_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9415_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Y11_9490_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9415_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9415_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9512_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9527_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Z0x2_9532_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Z0x2_9532_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Z1_9522_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Z1_9522_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9424_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9424_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9424_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9424_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9420_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9420_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9420_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9420_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS08_9418_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS08_9418_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS08_9418_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS08_9418_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Y00x2_9500_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9507_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9512_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS09_9419_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS09_9419_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS09_9419_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS09_9419_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Y00x2_9500_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9507_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9512_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9512_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9512_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9420_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9420_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Y11_9490_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9420_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9420_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9420_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9420_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9492_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9420_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9420_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Y12x2_9511_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Z1_9522_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Z0x2_9532_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Z0x2_9532_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Z1_9522_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9524_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9423_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9423_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9423_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9423_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS10_9421_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS10_9421_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS10_9421_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS10_9421_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9502_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9507_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Y12x2_9511_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Y12x2_9511_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS11_9422_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS11_9422_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS11_9422_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS11_9422_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9502_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9507_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Y12x2_9511_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Y02x2_9510_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Y02x2_9510_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Y02x2_9510_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9423_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9423_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9492_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9423_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9423_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9423_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9423_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9492_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9423_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9423_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Y02x2_9510_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9524_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9534_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9534_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9524_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9524_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Z0_9519_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Z0_9519_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9424_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9424_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9492_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9424_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9424_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9424_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9424_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Y10_9487_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9424_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9424_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9512_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Z0_9519_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9534_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9534_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Z0_9519_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9521_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9433_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9433_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9433_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9433_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9429_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9429_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9429_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9429_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS12_9427_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS12_9427_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS12_9427_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS12_9427_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9502_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9502_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9512_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9512_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS13_9428_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS13_9428_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS13_9428_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS13_9428_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9502_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9502_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9512_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9507_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9507_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9507_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9429_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9429_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Y10_9487_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9429_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9429_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9429_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9429_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Y10_9487_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9429_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9429_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9507_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9521_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Z3_9528_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Z3_9528_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9521_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9521_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9432_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9432_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9432_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9432_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS14_9430_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS14_9430_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS14_9430_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS14_9430_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Y13_9496_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9502_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9507_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS15_9431_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS15_9431_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS15_9431_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS15_9431_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Y13_9496_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9502_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9507_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9507_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9507_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9432_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9432_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Y10_9487_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9432_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9432_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9432_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9432_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9489_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9432_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9432_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Y11x2_9506_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9517_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Z3_9528_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Z3_9528_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9517_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9517_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9517_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9433_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9433_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9489_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9433_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9433_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9433_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9433_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9489_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9433_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9433_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Y11x2_9506_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9517_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9534_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9534_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9517_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9517_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9438_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9438_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9438_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9438_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS00x2_9436_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS00x2_9436_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS00x2_9436_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS00x2_9436_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9502_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Y11x2_9506_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Y11x2_9506_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9486_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS02x2_9437_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS02x2_9437_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS02x2_9437_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS02x2_9437_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9502_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9438_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9438_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9489_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9438_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9438_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9438_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9438_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Y03_9484_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9438_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9438_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9498_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9530_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9661_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Y12_9493_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9443_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9443_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9443_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9443_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS04x2_9441_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS04x2_9441_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS04x2_9441_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS04x2_9441_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Y10x2_9501_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS06x2_9442_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS06x2_9442_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS06x2_9442_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS06x2_9442_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS00x2_9623_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9634_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9443_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9443_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Y03_9484_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9443_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9443_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9443_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9443_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Y03_9484_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9443_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9443_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9502_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9448_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9448_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9448_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9448_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS08x2_9446_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS08x2_9446_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS08x2_9446_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS08x2_9446_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS10x2_9447_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS10x2_9447_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS10x2_9447_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS10x2_9447_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9448_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9448_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS04_9629_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9448_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9448_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9448_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9448_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS04_9629_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9448_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9448_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9630_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9661_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9630_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9624_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9453_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9453_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9453_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9453_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS12x2_9451_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS12x2_9451_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS12x2_9451_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9660_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9660_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS07x2_9658_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS07x2_9658_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS07x2_9658_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS07x2_9658_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS03_9755_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9634_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS14x2_9452_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS14x2_9452_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS14x2_9452_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS14x2_9452_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS00x2_9623_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9624_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9453_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9453_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS04_9629_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9453_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9453_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9453_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9453_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9453_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9453_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9657_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9652_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9652_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9458_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9458_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9458_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9458_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS01x2_9456_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS01x2_9456_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS01x2_9456_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS01x2_9456_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS00x2_9623_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9630_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS03x2_9457_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS03x2_9457_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS03x2_9457_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS03x2_9457_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9633_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9648_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9458_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9458_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9458_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9458_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9458_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9458_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9458_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9458_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9634_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9463_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9463_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9463_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9463_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS05x2_9461_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS05x2_9461_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS05x2_9461_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS05x2_9461_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9633_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9624_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS07x2_9462_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS07x2_9462_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS07x2_9462_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS07x2_9462_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9633_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9624_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9630_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9463_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9463_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9624_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9463_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9463_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9463_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9463_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9463_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9463_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9468_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9468_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9468_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9468_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS09x2_9466_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS09x2_9466_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS09x2_9466_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS09x2_9466_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS11x2_9467_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS11x2_9467_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS11x2_9467_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS11x2_9467_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9468_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9468_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9468_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9468_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9468_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9468_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9468_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9468_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9473_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9473_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9473_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9473_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS13x2_9471_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS13x2_9471_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS13x2_9471_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS13x2_9471_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS15x2_9472_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS15x2_9472_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS15x2_9472_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS15x2_9472_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9473_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9473_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9473_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9473_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9473_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9473_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9473_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9473_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9477_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9477_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9477_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9477_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Y00_9475_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Y00_9475_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9534_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9534_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9534_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9534_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9534_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9534_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9539_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9539_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9539_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9539_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Z1x2_9537_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Z1x2_9537_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Z1x2_9537_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Z1x2_9537_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Wc1_9538_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Wc1_9538_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Wc1_9538_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Wc1_9538_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9539_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9539_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9539_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9539_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9539_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9539_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9539_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9539_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9544_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9544_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9544_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9544_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Z2x2_9542_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Z2x2_9542_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Z2x2_9542_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Z2x2_9542_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Wc2_9543_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Wc2_9543_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Wc2_9543_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Wc2_9543_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9544_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9544_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9544_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9544_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9544_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9544_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9544_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9544_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9549_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9549_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9549_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9549_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Z3x2_9547_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Z3x2_9547_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Z3x2_9547_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Z3x2_9547_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Wc3_9548_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Wc3_9548_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Wc3_9548_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Wc3_9548_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9549_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9549_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9549_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9549_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9549_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9549_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9549_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9549_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9554_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9554_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9554_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9554_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_A0_9552_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_A0_9552_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_A0_9552_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_A0_9552_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Y00x2_9553_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Y00x2_9553_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Y00x2_9553_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Y00x2_9553_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9554_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9554_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9554_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9554_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9554_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9554_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9554_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9554_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9559_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9559_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9559_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9559_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_A1_9557_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_A1_9557_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_A1_9557_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_A1_9557_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Y01x2_9558_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Y01x2_9558_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Y01x2_9558_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Y01x2_9558_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9559_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9559_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9559_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9559_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9559_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9559_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9559_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9559_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9564_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9564_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9564_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9564_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_A2_9562_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_A2_9562_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_A2_9562_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_A2_9562_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Y02x2_9563_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Y02x2_9563_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Y02x2_9563_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Y02x2_9563_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9564_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9564_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9564_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9564_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9564_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9564_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9564_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9564_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9569_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9569_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9569_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9569_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_A3_9567_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_A3_9567_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_A3_9567_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_A3_9567_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Y03x2_9568_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Y03x2_9568_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Y03x2_9568_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Y03x2_9568_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9569_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9569_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9569_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9569_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9569_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9569_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9569_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9569_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9652_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9652_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9574_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9574_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9574_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9574_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_A0_9572_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_A0_9572_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_A0_9572_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_A0_9572_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS06_9647_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS06_9647_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Y10x2_9573_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Y10x2_9573_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Y10x2_9573_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Y10x2_9573_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9633_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9639_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS06_9647_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS06_9647_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_B01_9646_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_B01_9646_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9574_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9574_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS04_9629_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9574_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9574_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9574_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9574_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_B01_9628_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9574_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9574_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_B01_9646_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9657_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9657_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9652_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9652_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9579_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9579_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9579_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9579_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_A1_9577_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_A1_9577_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_A1_9577_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_A1_9577_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9633_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9639_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_B01_9646_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9648_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Y11x2_9578_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Y11x2_9578_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Y11x2_9578_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Y11x2_9578_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9633_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9643_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9648_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9648_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9648_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9652_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9579_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9579_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_B01_9628_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9579_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9579_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9579_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9579_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_B01_9628_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9579_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9579_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9652_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9652_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9657_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9657_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9652_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9584_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9584_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9584_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9584_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_A2_9582_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_A2_9582_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_A2_9582_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_A2_9582_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9633_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9643_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9652_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9652_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Y12x2_9583_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Y12x2_9583_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Y12x2_9583_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Y12x2_9583_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9643_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9643_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9643_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9643_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9643_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9584_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9584_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_B01_9628_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9584_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9584_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9584_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9584_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9630_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9584_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9584_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9651_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9657_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9657_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9651_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9651_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9589_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9589_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9589_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9589_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_A3_9587_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_A3_9587_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_A3_9587_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_A3_9587_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS05x2_9632_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9643_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9643_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9643_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Y13x2_9588_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Y13x2_9588_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Y13x2_9588_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Y13x2_9588_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS05x2_9632_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9634_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9643_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9643_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9642_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9589_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9589_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9630_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9589_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9589_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9589_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9589_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9630_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9589_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9589_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9642_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9651_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9657_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9657_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9651_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9598_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9598_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9598_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9598_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9594_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9594_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9594_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9594_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_B00_9592_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_B00_9592_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_B00_9592_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_B00_9592_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS05x2_9632_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9661_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9642_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9642_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS00_9593_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS00_9593_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS00_9593_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS00_9593_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9634_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9642_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9642_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9642_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9594_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9594_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9630_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9594_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9594_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9594_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9594_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9634_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9594_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9594_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9642_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9651_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS07_9656_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS07_9656_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9651_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9651_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9597_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9597_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9597_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9597_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS00x2_9595_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS00x2_9595_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS00x2_9595_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS00x2_9595_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS05x2_9632_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9634_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS06x2_9641_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS01x2_9596_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS01x2_9596_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS01x2_9596_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS01x2_9596_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS04x2_9631_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS06x2_9641_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS06x2_9641_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS06x2_9641_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS05x2_9640_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS05x2_9640_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9597_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9597_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9634_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9597_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9597_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9597_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9597_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9634_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9597_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9597_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS05x2_9640_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS07_9656_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS07_9656_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS07x2_9650_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS07x2_9650_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS07x2_9650_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS07x2_9650_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9598_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9598_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9634_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9598_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9598_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9598_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9598_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9625_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9598_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9598_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS05x2_9640_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS06x2_9649_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_B11_9655_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IMX03_9756_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS06x2_9649_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS06x2_9649_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9607_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9607_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9607_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9607_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9603_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9603_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9603_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9603_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_B10_9601_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_B10_9601_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_B10_9601_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_B10_9601_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS04x2_9631_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9642_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9642_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9642_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS01_9602_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS01_9602_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS01_9602_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS01_9602_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9634_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9642_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9639_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9639_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9639_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9603_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9603_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9625_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9603_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9603_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9603_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9603_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9625_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9603_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9603_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9639_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS06x2_9649_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_B11_9655_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_B11_9655_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9651_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9651_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9606_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9606_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9606_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9606_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS01x2_9604_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS01x2_9604_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS01x2_9604_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS01x2_9604_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS04x2_9631_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9639_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS02x2_9605_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS02x2_9605_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS02x2_9605_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS02x2_9605_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS04x2_9631_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9639_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9639_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9639_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS05_9638_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9606_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9606_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9625_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9606_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9606_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9606_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9606_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9625_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9606_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9606_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS05_9638_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9651_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9657_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_B11_9655_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9651_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9648_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9648_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9648_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9607_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9607_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9625_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9607_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9607_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9607_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9607_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9625_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9607_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9607_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS05_9638_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9648_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9657_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9657_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9648_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9616_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9616_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9616_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9616_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9612_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9612_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9612_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9612_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_B00_9610_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_B00_9610_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_B00_9610_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_B00_9610_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9633_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9634_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS05_9638_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_B11_9637_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS02_9611_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS02_9611_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS02_9611_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS02_9611_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9633_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_B11_9637_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_B11_9637_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_B11_9637_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9639_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9612_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9612_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9625_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9612_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9612_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9612_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9612_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9624_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9612_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9612_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9639_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9648_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9660_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9660_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9648_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9633_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9615_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9615_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9615_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9615_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS02x2_9613_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS02x2_9613_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS02x2_9613_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS02x2_9613_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9633_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS03x2_9614_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS03x2_9614_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS03x2_9614_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS03x2_9614_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9633_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9615_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9615_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9624_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9615_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9615_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9615_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9615_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9624_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9615_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9615_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9630_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9661_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS03_9755_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9630_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9630_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_l_round_9772_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9616_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9616_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9616_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9616_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9616_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9616_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9616_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9616_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9769_complete/ack
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IMX06_9774_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IMX04_9762_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9625_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9625_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9625_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9625_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9621_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9621_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9621_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9621_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_B10_9619_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_B10_9619_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_B10_9619_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_B10_9619_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9775_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS03_9755_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS03_9620_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS03_9620_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS03_9620_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS03_9620_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS05_9767_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9621_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9621_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9621_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9621_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9621_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9621_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9621_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9621_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9624_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9624_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9624_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9624_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS03x2_9622_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS03x2_9622_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS03x2_9622_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS03x2_9622_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS00x2_9623_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS04x2_9659_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS04x2_9659_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS04x2_9659_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS04x2_9659_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9660_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9660_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9660_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9660_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9660_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9660_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9660_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9660_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9661_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9661_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9661_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9661_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9661_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9661_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9661_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9661_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9670_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9670_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9670_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9670_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9666_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9666_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9666_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9666_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_B02_9664_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_B02_9664_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_B02_9664_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_B02_9664_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS08_9665_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS08_9665_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS08_9665_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS08_9665_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9666_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9666_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9666_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9666_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9666_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9666_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9666_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9666_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9669_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9669_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9669_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9669_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS08x2_9667_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS08x2_9667_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS08x2_9667_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS08x2_9667_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS09x2_9668_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS09x2_9668_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS09x2_9668_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS09x2_9668_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9669_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9669_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9669_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9669_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9669_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9669_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9669_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9669_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9670_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9670_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9670_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9670_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9670_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9670_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9670_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9670_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9679_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9679_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9679_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9679_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9675_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9675_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9675_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9675_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_B12_9673_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_B12_9673_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_B12_9673_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_B12_9673_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS09_9674_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS09_9674_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS09_9674_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS09_9674_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9675_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9675_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9675_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9675_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9675_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9675_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9675_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9675_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9678_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9678_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9678_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9678_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS09x2_9676_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS09x2_9676_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS09x2_9676_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS09x2_9676_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS10x2_9677_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS10x2_9677_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS10x2_9677_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS10x2_9677_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9678_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9678_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9678_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9678_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9678_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9678_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9678_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9678_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9679_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9679_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9679_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9679_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9679_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9679_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9679_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9679_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9688_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9688_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9688_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9688_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9684_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9684_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9684_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9684_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_B02_9682_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_B02_9682_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_B02_9682_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_B02_9682_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS10_9683_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS10_9683_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS10_9683_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS10_9683_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9684_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9684_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9684_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9684_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9684_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9684_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9684_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9684_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9687_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9687_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9687_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9687_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS10x2_9685_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS10x2_9685_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS10x2_9685_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS10x2_9685_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS11x2_9686_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS11x2_9686_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS11x2_9686_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS11x2_9686_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9687_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9687_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9687_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9687_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9687_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9687_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9687_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9687_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9688_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9688_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9688_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9688_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9688_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9688_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9688_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9688_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9697_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9697_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9697_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9697_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9693_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9693_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9693_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9693_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_B12_9691_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_B12_9691_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_B12_9691_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_B12_9691_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS11_9692_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS11_9692_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS11_9692_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS11_9692_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9763_start/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IMX05_9768_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9769_complete/req
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9769_complete/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9769_complete/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9693_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9693_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_l_round_9760_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9693_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9693_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9693_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9693_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9763_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9693_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9693_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9769_start/ack
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_l_round_9772_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IMX06_9774_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IMX06_9774_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_l_round_9772_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_l_round_9772_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9696_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9696_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9696_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9696_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS11x2_9694_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS11x2_9694_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS11x2_9694_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS11x2_9694_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS05_9767_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS05_9767_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9769_start/req
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9769_start/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS08x2_9695_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS08x2_9695_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS08x2_9695_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS08x2_9695_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_l_round_9766_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS05_9767_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9769_start/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IMX05_9768_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IMX05_9768_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9696_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9696_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9763_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9696_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9696_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9696_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9696_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9763_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9696_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9696_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IMX05_9768_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9775_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9775_start/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9775_start/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9775_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9775_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_l_round_9766_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_l_round_9766_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9697_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9697_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9763_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9697_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9697_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9697_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9697_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9757_complete/ack
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9697_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9697_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IMX04_9762_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IMX06_9774_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISX0_9916_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IMX04_9762_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_l_round_9766_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9706_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9706_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9706_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9706_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9702_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9702_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9702_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9702_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_B03_9700_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_B03_9700_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_B03_9700_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_B03_9700_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9769_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS12_9701_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS12_9701_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS12_9701_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS12_9701_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9702_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9702_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9757_complete/req
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9702_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9702_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9702_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9702_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9757_complete/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9702_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9702_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IMX04_9762_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS06_9773_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS04_9761_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9769_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9705_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9705_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9705_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9705_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS12x2_9703_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS12x2_9703_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS12x2_9703_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS12x2_9703_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9769_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS13x2_9704_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS13x2_9704_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS13x2_9704_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS13x2_9704_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9769_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9705_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9705_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9757_complete/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9705_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9705_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9705_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9705_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9757_start/ack
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9705_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9705_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS04_9761_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS06_9773_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS04_9761_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9763_complete/ack
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9763_complete/req
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9763_complete/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9706_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9706_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9757_start/req
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9706_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9706_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9706_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9706_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9757_start/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9706_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9706_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS04_9761_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS06_9773_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_l_round_9760_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9763_complete/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9715_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9715_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9715_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9715_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9711_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9711_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9711_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9711_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_B13_9709_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_B13_9709_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_B13_9709_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_B13_9709_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS13_9710_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS13_9710_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS13_9710_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS13_9710_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9711_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9711_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9757_start/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9711_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9711_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9711_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9711_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IMX03_9756_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9711_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9711_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_l_round_9760_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS06_9773_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u16_u32_9913_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_l_round_9760_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9763_start/ack
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9714_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9714_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9714_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9714_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS13x2_9712_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS13x2_9712_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS13x2_9712_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS13x2_9712_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9763_start/req
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS14x2_9713_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS14x2_9713_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS14x2_9713_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS14x2_9713_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9763_start/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9714_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9714_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IMX03_9756_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9714_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9714_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9714_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9714_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IMX03_9756_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9714_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9714_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u16_u32_9913_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u64_u128_9922_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9715_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9715_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9715_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9715_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9715_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9715_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISX0_9916_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9715_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9715_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISX0_9916_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9724_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9724_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9724_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9724_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9720_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9720_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9720_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9720_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_B03_9718_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_B03_9718_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_B03_9718_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_B03_9718_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u32_u64_9918_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS14_9719_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS14_9719_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS14_9719_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS14_9719_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u64_u128_9922_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u32_u64_9918_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9720_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9720_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9720_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9720_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9720_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9720_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9720_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9720_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u8_u16_9912_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9723_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9723_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9723_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9723_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS14x2_9721_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS14x2_9721_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS14x2_9721_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS14x2_9721_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u32_u64_9918_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u16_u32_9913_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS15x2_9722_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS15x2_9722_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS15x2_9722_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS15x2_9722_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9723_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9723_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9723_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9723_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9723_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9723_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9723_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9723_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u32_u64_9921_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u32_u64_9918_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9724_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9724_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9724_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9724_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9724_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9724_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9724_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9724_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9733_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9733_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9733_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9733_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9729_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9729_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9729_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9729_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_B13_9727_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_B13_9727_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_B13_9727_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_B13_9727_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS15_9728_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS15_9728_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS15_9728_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS15_9728_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u32_u64_9921_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u128_u128_9927_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u16_u32_9913_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u16_u32_9913_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9729_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9729_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u8_u16_9912_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9729_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9729_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9729_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9729_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u16_u32_9913_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9729_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9729_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u16_u32_9913_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u32_u64_9921_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9732_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9732_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9732_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9732_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS15x2_9730_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS15x2_9730_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS15x2_9730_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS15x2_9730_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS12x2_9731_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS12x2_9731_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS12x2_9731_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS12x2_9731_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u32_u64_9921_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9732_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9732_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u64_u128_9922_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9732_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9732_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9732_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9732_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u64_u128_9922_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9732_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9732_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u16_u32_9913_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u128_u128_9927_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u32_u64_9921_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9733_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9733_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9733_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9733_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9733_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9733_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9733_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u8_u8_9733_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9739_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9739_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9739_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9739_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_l_round_9736_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_l_round_9736_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_l_round_9736_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_l_round_9736_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS00_9737_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS00_9737_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS00_9737_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS00_9737_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IMX00_9738_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IMX00_9738_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IMX00_9738_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IMX00_9738_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9739_start/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9739_start/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9739_start/req
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9739_start/ack
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9739_complete/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9739_complete/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9739_complete/req
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9739_complete/ack
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9745_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9745_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9745_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9745_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_l_round_9742_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_l_round_9742_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_l_round_9742_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_l_round_9742_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS01_9743_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS01_9743_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS01_9743_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS01_9743_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IMX01_9744_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IMX01_9744_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IMX01_9744_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IMX01_9744_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9745_start/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9745_start/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9745_start/req
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9745_start/ack
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9745_complete/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9745_complete/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9745_complete/req
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9745_complete/ack
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9751_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9751_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9751_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9751_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_l_round_9748_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_l_round_9748_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_l_round_9748_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_l_round_9748_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS02_9749_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS02_9749_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS02_9749_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS02_9749_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IMX02_9750_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IMX02_9750_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IMX02_9750_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IMX02_9750_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9751_start/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9751_start/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9751_start/req
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9751_start/ack
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9751_complete/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9751_complete/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9751_complete/req
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9751_complete/ack
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9757_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9757_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9757_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9757_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_l_round_9754_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_l_round_9754_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_l_round_9754_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_l_round_9754_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS03_9755_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9775_start/req
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9775_start/ack
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9775_complete/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9775_complete/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9775_complete/req
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9775_complete/ack
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9781_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9781_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9781_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9781_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_l_round_9778_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_l_round_9778_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_l_round_9778_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_l_round_9778_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS07_9779_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS07_9779_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS07_9779_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS07_9779_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IMX07_9780_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IMX07_9780_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IMX07_9780_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IMX07_9780_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9781_start/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9781_start/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9781_start/req
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9781_start/ack
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9781_complete/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9781_complete/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9781_complete/req
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9781_complete/ack
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9787_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9787_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9787_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9787_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_l_round_9784_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_l_round_9784_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_l_round_9784_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_l_round_9784_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS08_9785_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS08_9785_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS08_9785_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS08_9785_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IMX08_9786_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IMX08_9786_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IMX08_9786_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IMX08_9786_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9787_start/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9787_start/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9787_start/req
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9787_start/ack
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9787_complete/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9787_complete/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9787_complete/req
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9787_complete/ack
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9793_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9793_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9793_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9793_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_l_round_9790_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_l_round_9790_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_l_round_9790_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_l_round_9790_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS09_9791_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS09_9791_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS09_9791_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS09_9791_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IMX09_9792_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IMX09_9792_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IMX09_9792_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IMX09_9792_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9793_start/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9793_start/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9793_start/req
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9793_start/ack
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9793_complete/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9793_complete/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9793_complete/req
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9793_complete/ack
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9799_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9799_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9799_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9799_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_l_round_9796_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_l_round_9796_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_l_round_9796_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_l_round_9796_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS10_9797_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS10_9797_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS10_9797_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS10_9797_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IMX10_9798_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IMX10_9798_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IMX10_9798_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IMX10_9798_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9799_start/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9799_start/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9799_start/req
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9799_start/ack
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9799_complete/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9799_complete/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9799_complete/req
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9799_complete/ack
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9805_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9805_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9805_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9805_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_l_round_9802_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_l_round_9802_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_l_round_9802_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_l_round_9802_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS11_9803_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS11_9803_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS11_9803_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS11_9803_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IMX11_9804_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IMX11_9804_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IMX11_9804_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IMX11_9804_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9805_start/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9805_start/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9805_start/req
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9805_start/ack
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9805_complete/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9805_complete/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9805_complete/req
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9805_complete/ack
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9811_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9811_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9811_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9811_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_l_round_9808_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_l_round_9808_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_l_round_9808_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_l_round_9808_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS12_9809_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS12_9809_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS12_9809_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS12_9809_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IMX12_9810_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IMX12_9810_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IMX12_9810_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IMX12_9810_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9811_start/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9811_start/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9811_start/req
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9811_start/ack
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9811_complete/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9811_complete/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9811_complete/req
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9811_complete/ack
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9817_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9817_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9817_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9817_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_l_round_9814_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_l_round_9814_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_l_round_9814_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_l_round_9814_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS13_9815_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS13_9815_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS13_9815_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS13_9815_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IMX13_9816_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IMX13_9816_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IMX13_9816_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IMX13_9816_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9817_start/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9817_start/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9817_start/req
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9817_start/ack
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9817_complete/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9817_complete/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9817_complete/req
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9817_complete/ack
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9823_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9823_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9823_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9823_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_l_round_9820_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_l_round_9820_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_l_round_9820_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_l_round_9820_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS14_9821_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS14_9821_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS14_9821_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS14_9821_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IMX14_9822_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IMX14_9822_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IMX14_9822_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IMX14_9822_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9823_start/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9823_start/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9823_start/req
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9823_start/ack
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9823_complete/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9823_complete/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9823_complete/req
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9823_complete/ack
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9829_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9829_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9829_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9829_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_l_round_9826_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_l_round_9826_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_l_round_9826_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_l_round_9826_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS15_9827_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS15_9827_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS15_9827_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IS15_9827_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IMX15_9828_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IMX15_9828_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IMX15_9828_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_IMX15_9828_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9829_start/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9829_start/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9829_start/req
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9829_start/ack
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9829_complete/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9829_complete/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9829_complete/req
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/MUX_9829_complete/ack
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9833_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9833_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9833_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9833_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISbox_in00_9831_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISbox_in00_9831_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISbox_in00_9831_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISbox_in00_9831_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9836_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9836_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9836_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9836_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISbox_in01_9834_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISbox_in01_9834_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISbox_in01_9834_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISbox_in01_9834_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9839_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9839_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9839_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9839_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISbox_in02_9837_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISbox_in02_9837_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISbox_in02_9837_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISbox_in02_9837_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9842_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9842_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9842_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9842_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u128_u128_9927_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u32_u64_9921_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISbox_in03_9840_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISbox_in03_9840_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISbox_in03_9840_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISbox_in03_9840_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u32_u64_9921_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISX3_9920_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u128_u128_9927_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9845_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9845_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9845_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9845_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISX3_9920_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISbox_in04_9843_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISbox_in04_9843_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISbox_in04_9843_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISbox_in04_9843_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISX3_9920_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_key_in_9926_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISX3_9920_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_key_in_9926_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9848_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9848_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9848_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9848_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_key_in_9926_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISX2_9919_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISbox_in05_9846_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISbox_in05_9846_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISbox_in05_9846_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISbox_in05_9846_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISX2_9919_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_key_in_9926_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISX2_9919_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_OUT_9925_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9851_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9851_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9851_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9851_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_OUT_9925_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISX2_9919_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISbox_in06_9849_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISbox_in06_9849_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISbox_in06_9849_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISbox_in06_9849_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u32_u64_9921_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_OUT_9925_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u32_u64_9921_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_OUT_9925_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9854_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9854_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9854_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9854_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u32_u64_9921_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISbox_in07_9852_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISbox_in07_9852_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISbox_in07_9852_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISbox_in07_9852_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u32_u64_9921_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u128_u128_9927_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u32_u64_9918_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9857_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9857_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9857_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9857_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u128_u128_9927_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u32_u64_9918_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISbox_in08_9855_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISbox_in08_9855_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISbox_in08_9855_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISbox_in08_9855_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u32_u64_9918_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u64_u128_9922_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u32_u64_9918_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u64_u128_9922_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9860_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9860_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9860_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9860_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u64_u128_9922_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u32_u64_9918_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISbox_in09_9858_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISbox_in09_9858_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISbox_in09_9858_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISbox_in09_9858_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u32_u64_9918_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u64_u128_9922_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u32_u64_9918_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9863_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9863_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9863_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9863_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u64_u128_9922_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u32_u64_9918_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISbox_in10_9861_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISbox_in10_9861_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISbox_in10_9861_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISbox_in10_9861_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISX1_9917_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u64_u128_9922_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISX1_9917_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u64_u128_9922_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9866_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9866_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9866_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9866_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u64_u128_9922_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISX1_9917_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISbox_in11_9864_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISbox_in11_9864_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISbox_in11_9864_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISbox_in11_9864_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISX1_9917_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISX0_9916_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u32_u64_9921_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9869_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9869_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9869_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9869_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISbox_in12_9867_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISbox_in12_9867_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISbox_in12_9867_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISbox_in12_9867_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9872_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9872_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9872_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9872_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISbox_in13_9870_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISbox_in13_9870_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISbox_in13_9870_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISbox_in13_9870_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9875_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9875_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9875_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9875_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISbox_in14_9873_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISbox_in14_9873_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISbox_in14_9873_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISbox_in14_9873_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9878_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9878_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9878_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/call_stmt_9878_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISbox_in15_9876_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISbox_in15_9876_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISbox_in15_9876_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_ISbox_in15_9876_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u16_u32_9886_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u16_u32_9886_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u16_u32_9886_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u16_u32_9886_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u8_u16_9882_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u8_u16_9882_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u8_u16_9882_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u8_u16_9882_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Sout00_9880_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Sout00_9880_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Sout00_9880_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Sout00_9880_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Sout01_9881_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Sout01_9881_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Sout01_9881_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Sout01_9881_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u8_u16_9882_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u8_u16_9882_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u8_u16_9882_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u8_u16_9882_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u8_u16_9882_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u8_u16_9882_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u8_u16_9882_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u8_u16_9882_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u8_u16_9885_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u8_u16_9885_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u8_u16_9885_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u8_u16_9885_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Sout02_9883_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Sout02_9883_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Sout02_9883_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Sout02_9883_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Sout03_9884_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Sout03_9884_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Sout03_9884_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Sout03_9884_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u8_u16_9885_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u8_u16_9885_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u8_u16_9885_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u8_u16_9885_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u8_u16_9885_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u8_u16_9885_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u8_u16_9885_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u8_u16_9885_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u16_u32_9886_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u16_u32_9886_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u16_u32_9886_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u16_u32_9886_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u16_u32_9886_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u16_u32_9886_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u16_u32_9886_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u16_u32_9886_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u16_u32_9895_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u16_u32_9895_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u16_u32_9895_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u16_u32_9895_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u8_u16_9891_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u8_u16_9891_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u8_u16_9891_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u8_u16_9891_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Sout04_9889_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Sout04_9889_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Sout04_9889_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Sout04_9889_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Sout05_9890_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Sout05_9890_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Sout05_9890_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Sout05_9890_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u8_u16_9891_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u8_u16_9891_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u8_u16_9891_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u8_u16_9891_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u8_u16_9891_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u8_u16_9891_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u8_u16_9891_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u8_u16_9891_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u8_u16_9894_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u8_u16_9894_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u8_u16_9894_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u8_u16_9894_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Sout06_9892_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Sout06_9892_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Sout06_9892_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Sout06_9892_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Sout07_9893_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Sout07_9893_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Sout07_9893_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Sout07_9893_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u8_u16_9894_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u8_u16_9894_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u8_u16_9894_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u8_u16_9894_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u8_u16_9894_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u8_u16_9894_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u8_u16_9894_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u8_u16_9894_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u16_u32_9895_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u16_u32_9895_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u16_u32_9895_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u16_u32_9895_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u16_u32_9895_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u16_u32_9895_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u16_u32_9895_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u16_u32_9895_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u16_u32_9904_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u16_u32_9904_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u16_u32_9904_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u16_u32_9904_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u8_u16_9900_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u8_u16_9900_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u8_u16_9900_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u8_u16_9900_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Sout08_9898_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Sout08_9898_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Sout08_9898_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Sout08_9898_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Sout09_9899_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Sout09_9899_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Sout09_9899_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Sout09_9899_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u8_u16_9900_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u8_u16_9900_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u8_u16_9900_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u8_u16_9900_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u8_u16_9900_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u8_u16_9900_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u8_u16_9900_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u8_u16_9900_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u8_u16_9903_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u8_u16_9903_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u8_u16_9903_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u8_u16_9903_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Sout10_9901_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Sout10_9901_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Sout10_9901_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Sout10_9901_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Sout11_9902_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Sout11_9902_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Sout11_9902_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Sout11_9902_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u8_u16_9903_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u8_u16_9903_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u8_u16_9903_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u8_u16_9903_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u8_u16_9903_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u8_u16_9903_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u8_u16_9903_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u8_u16_9903_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u16_u32_9904_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u16_u32_9904_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u16_u32_9904_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u16_u32_9904_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u16_u32_9904_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u16_u32_9904_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u16_u32_9904_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u16_u32_9904_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u16_u32_9913_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u16_u32_9913_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u16_u32_9913_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u16_u32_9913_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u8_u16_9909_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u8_u16_9909_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u8_u16_9909_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u8_u16_9909_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Sout12_9907_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Sout12_9907_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Sout12_9907_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Sout12_9907_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Sout13_9908_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Sout13_9908_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Sout13_9908_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Sout13_9908_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u8_u16_9909_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u8_u16_9909_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u8_u16_9909_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u8_u16_9909_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u8_u16_9909_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u8_u16_9909_Update/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u8_u16_9909_Update/cr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u8_u16_9909_Update/ca
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u8_u16_9912_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u8_u16_9912_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u8_u16_9912_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u8_u16_9912_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Sout14_9910_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Sout14_9910_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Sout14_9910_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Sout14_9910_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Sout15_9911_sample_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Sout15_9911_sample_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Sout15_9911_update_start_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/R_Sout15_9911_update_completed_
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u8_u16_9912_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u8_u16_9912_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u8_u16_9912_Sample/rr
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u8_u16_9912_Sample/ra
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u8_u16_9912_Update/$entry
      -- CP-element group 0: 	 assign_stmt_9274_to_assign_stmt_9928/CONCAT_u8_u16_9912_Update/$exit
      -- 
    -- logger for CP element group dec_round_CP_192_elements(0)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and dec_round_CP_192_elements(0)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:dec_round:CP:dec_round_CP_192_elements(0) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:dec_round:CP:XOR_u128_u128_9927_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:dec_round:CP:XOR_u128_u128_9927_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    cr_3324_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => dec_round_CP_192_elements(0), ack => XOR_u128_u128_9927_inst_req_1); -- 
    rr_3319_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => dec_round_CP_192_elements(0), ack => XOR_u128_u128_9927_inst_req_0); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u128_u128_9927_Sample/ra
      -- CP-element group 1: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u128_u128_9927_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u128_u128_9927_sample_completed_
      -- 
    -- logger for CP element group dec_round_CP_192_elements(1)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and dec_round_CP_192_elements(1)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:dec_round:CP:dec_round_CP_192_elements(1) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:dec_round:CP:XOR_u128_u128_9927_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_3320_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => XOR_u128_u128_9927_inst_ack_0, ack => dec_round_CP_192_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2:  members (5) 
      -- CP-element group 2: 	 $exit
      -- CP-element group 2: 	 assign_stmt_9274_to_assign_stmt_9928/$exit
      -- CP-element group 2: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u128_u128_9927_Update/ca
      -- CP-element group 2: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u128_u128_9927_Update/$exit
      -- CP-element group 2: 	 assign_stmt_9274_to_assign_stmt_9928/XOR_u128_u128_9927_update_completed_
      -- 
    -- logger for CP element group dec_round_CP_192_elements(2)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and dec_round_CP_192_elements(2)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:dec_round:CP:dec_round_CP_192_elements(2) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:dec_round:CP:XOR_u128_u128_9927_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_3325_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => XOR_u128_u128_9927_inst_ack_1, ack => dec_round_CP_192_elements(2)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal A0_9535 : std_logic_vector(7 downto 0);
    signal A1_9540 : std_logic_vector(7 downto 0);
    signal A2_9545 : std_logic_vector(7 downto 0);
    signal A3_9550 : std_logic_vector(7 downto 0);
    signal B00_9555 : std_logic_vector(7 downto 0);
    signal B01_9560 : std_logic_vector(7 downto 0);
    signal B02_9565 : std_logic_vector(7 downto 0);
    signal B03_9570 : std_logic_vector(7 downto 0);
    signal B10_9575 : std_logic_vector(7 downto 0);
    signal B11_9580 : std_logic_vector(7 downto 0);
    signal B12_9585 : std_logic_vector(7 downto 0);
    signal B13_9590 : std_logic_vector(7 downto 0);
    signal CONCAT_u32_u64_9918_wire : std_logic_vector(63 downto 0);
    signal CONCAT_u32_u64_9921_wire : std_logic_vector(63 downto 0);
    signal CONCAT_u8_u16_9882_wire : std_logic_vector(15 downto 0);
    signal CONCAT_u8_u16_9885_wire : std_logic_vector(15 downto 0);
    signal CONCAT_u8_u16_9891_wire : std_logic_vector(15 downto 0);
    signal CONCAT_u8_u16_9894_wire : std_logic_vector(15 downto 0);
    signal CONCAT_u8_u16_9900_wire : std_logic_vector(15 downto 0);
    signal CONCAT_u8_u16_9903_wire : std_logic_vector(15 downto 0);
    signal CONCAT_u8_u16_9909_wire : std_logic_vector(15 downto 0);
    signal CONCAT_u8_u16_9912_wire : std_logic_vector(15 downto 0);
    signal IMX00_9599 : std_logic_vector(7 downto 0);
    signal IMX01_9608 : std_logic_vector(7 downto 0);
    signal IMX02_9617 : std_logic_vector(7 downto 0);
    signal IMX03_9626 : std_logic_vector(7 downto 0);
    signal IMX04_9635 : std_logic_vector(7 downto 0);
    signal IMX05_9644 : std_logic_vector(7 downto 0);
    signal IMX06_9653 : std_logic_vector(7 downto 0);
    signal IMX07_9662 : std_logic_vector(7 downto 0);
    signal IMX08_9671 : std_logic_vector(7 downto 0);
    signal IMX09_9680 : std_logic_vector(7 downto 0);
    signal IMX10_9689 : std_logic_vector(7 downto 0);
    signal IMX11_9698 : std_logic_vector(7 downto 0);
    signal IMX12_9707 : std_logic_vector(7 downto 0);
    signal IMX13_9716 : std_logic_vector(7 downto 0);
    signal IMX14_9725 : std_logic_vector(7 downto 0);
    signal IMX15_9734 : std_logic_vector(7 downto 0);
    signal IS00_9290 : std_logic_vector(7 downto 0);
    signal IS00x2_9353 : std_logic_vector(7 downto 0);
    signal IS01_9294 : std_logic_vector(7 downto 0);
    signal IS01x2_9356 : std_logic_vector(7 downto 0);
    signal IS02_9298 : std_logic_vector(7 downto 0);
    signal IS02x2_9359 : std_logic_vector(7 downto 0);
    signal IS03_9302 : std_logic_vector(7 downto 0);
    signal IS03x2_9362 : std_logic_vector(7 downto 0);
    signal IS04_9306 : std_logic_vector(7 downto 0);
    signal IS04x2_9365 : std_logic_vector(7 downto 0);
    signal IS05_9310 : std_logic_vector(7 downto 0);
    signal IS05x2_9368 : std_logic_vector(7 downto 0);
    signal IS06_9314 : std_logic_vector(7 downto 0);
    signal IS06x2_9371 : std_logic_vector(7 downto 0);
    signal IS07_9318 : std_logic_vector(7 downto 0);
    signal IS07x2_9374 : std_logic_vector(7 downto 0);
    signal IS08_9322 : std_logic_vector(7 downto 0);
    signal IS08x2_9377 : std_logic_vector(7 downto 0);
    signal IS09_9326 : std_logic_vector(7 downto 0);
    signal IS09x2_9380 : std_logic_vector(7 downto 0);
    signal IS10_9330 : std_logic_vector(7 downto 0);
    signal IS10x2_9383 : std_logic_vector(7 downto 0);
    signal IS11_9334 : std_logic_vector(7 downto 0);
    signal IS11x2_9386 : std_logic_vector(7 downto 0);
    signal IS12_9338 : std_logic_vector(7 downto 0);
    signal IS12x2_9389 : std_logic_vector(7 downto 0);
    signal IS13_9342 : std_logic_vector(7 downto 0);
    signal IS13x2_9392 : std_logic_vector(7 downto 0);
    signal IS14_9346 : std_logic_vector(7 downto 0);
    signal IS14x2_9395 : std_logic_vector(7 downto 0);
    signal IS15_9350 : std_logic_vector(7 downto 0);
    signal IS15x2_9398 : std_logic_vector(7 downto 0);
    signal ISX0_9887 : std_logic_vector(31 downto 0);
    signal ISX1_9896 : std_logic_vector(31 downto 0);
    signal ISX2_9905 : std_logic_vector(31 downto 0);
    signal ISX3_9914 : std_logic_vector(31 downto 0);
    signal ISa_9274 : std_logic_vector(31 downto 0);
    signal ISb_9278 : std_logic_vector(31 downto 0);
    signal ISbox_in00_9740 : std_logic_vector(7 downto 0);
    signal ISbox_in01_9746 : std_logic_vector(7 downto 0);
    signal ISbox_in02_9752 : std_logic_vector(7 downto 0);
    signal ISbox_in03_9758 : std_logic_vector(7 downto 0);
    signal ISbox_in04_9764 : std_logic_vector(7 downto 0);
    signal ISbox_in05_9770 : std_logic_vector(7 downto 0);
    signal ISbox_in06_9776 : std_logic_vector(7 downto 0);
    signal ISbox_in07_9782 : std_logic_vector(7 downto 0);
    signal ISbox_in08_9788 : std_logic_vector(7 downto 0);
    signal ISbox_in09_9794 : std_logic_vector(7 downto 0);
    signal ISbox_in10_9800 : std_logic_vector(7 downto 0);
    signal ISbox_in11_9806 : std_logic_vector(7 downto 0);
    signal ISbox_in12_9812 : std_logic_vector(7 downto 0);
    signal ISbox_in13_9818 : std_logic_vector(7 downto 0);
    signal ISbox_in14_9824 : std_logic_vector(7 downto 0);
    signal ISbox_in15_9830 : std_logic_vector(7 downto 0);
    signal ISc_9282 : std_logic_vector(31 downto 0);
    signal ISd_9286 : std_logic_vector(31 downto 0);
    signal OUT_9923 : std_logic_vector(127 downto 0);
    signal Sout00_9833 : std_logic_vector(7 downto 0);
    signal Sout01_9872 : std_logic_vector(7 downto 0);
    signal Sout02_9863 : std_logic_vector(7 downto 0);
    signal Sout03_9854 : std_logic_vector(7 downto 0);
    signal Sout04_9845 : std_logic_vector(7 downto 0);
    signal Sout05_9836 : std_logic_vector(7 downto 0);
    signal Sout06_9875 : std_logic_vector(7 downto 0);
    signal Sout07_9866 : std_logic_vector(7 downto 0);
    signal Sout08_9857 : std_logic_vector(7 downto 0);
    signal Sout09_9848 : std_logic_vector(7 downto 0);
    signal Sout10_9839 : std_logic_vector(7 downto 0);
    signal Sout11_9878 : std_logic_vector(7 downto 0);
    signal Sout12_9869 : std_logic_vector(7 downto 0);
    signal Sout13_9860 : std_logic_vector(7 downto 0);
    signal Sout14_9851 : std_logic_vector(7 downto 0);
    signal Sout15_9842 : std_logic_vector(7 downto 0);
    signal Wc0_9407 : std_logic_vector(7 downto 0);
    signal Wc1_9416 : std_logic_vector(7 downto 0);
    signal Wc2_9425 : std_logic_vector(7 downto 0);
    signal Wc3_9434 : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_9402_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_9405_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_9411_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_9414_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_9420_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_9423_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_9429_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_9432_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_9594_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_9597_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_9603_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_9606_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_9612_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_9615_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_9621_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_9624_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_9630_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_9633_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_9639_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_9642_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_9648_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_9651_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_9657_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_9660_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_9666_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_9669_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_9675_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_9678_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_9684_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_9687_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_9693_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_9696_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_9702_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_9705_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_9711_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_9714_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_9720_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_9723_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_9729_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_9732_wire : std_logic_vector(7 downto 0);
    signal Y00_9439 : std_logic_vector(7 downto 0);
    signal Y00x2_9477 : std_logic_vector(7 downto 0);
    signal Y01_9444 : std_logic_vector(7 downto 0);
    signal Y01x2_9480 : std_logic_vector(7 downto 0);
    signal Y02_9449 : std_logic_vector(7 downto 0);
    signal Y02x2_9483 : std_logic_vector(7 downto 0);
    signal Y03_9454 : std_logic_vector(7 downto 0);
    signal Y03x2_9486 : std_logic_vector(7 downto 0);
    signal Y10_9459 : std_logic_vector(7 downto 0);
    signal Y10x2_9489 : std_logic_vector(7 downto 0);
    signal Y11_9464 : std_logic_vector(7 downto 0);
    signal Y11x2_9492 : std_logic_vector(7 downto 0);
    signal Y12_9469 : std_logic_vector(7 downto 0);
    signal Y12x2_9495 : std_logic_vector(7 downto 0);
    signal Y13_9474 : std_logic_vector(7 downto 0);
    signal Y13x2_9498 : std_logic_vector(7 downto 0);
    signal Z0_9503 : std_logic_vector(7 downto 0);
    signal Z0x2_9521 : std_logic_vector(7 downto 0);
    signal Z1_9508 : std_logic_vector(7 downto 0);
    signal Z1x2_9524 : std_logic_vector(7 downto 0);
    signal Z2_9513 : std_logic_vector(7 downto 0);
    signal Z2x2_9527 : std_logic_vector(7 downto 0);
    signal Z3_9518 : std_logic_vector(7 downto 0);
    signal Z3x2_9530 : std_logic_vector(7 downto 0);
    signal xxdec_roundxxsel : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    xxdec_roundxxsel <= "01111111";
    -- logger for split-operator MUX_9739_inst flow-through 
    process(ISbox_in00_9740) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:MUX_9739_inst:flowthrough inputs: " & " l_round_buffer = "& Convert_SLV_To_Hex_String(l_round_buffer) & " IS00_9290 = "& Convert_SLV_To_Hex_String(IS00_9290) & " IMX00_9599 = "& Convert_SLV_To_Hex_String(IMX00_9599) & " outputs:" & " ISbox_in00_9740= "  & Convert_SLV_To_Hex_String(ISbox_in00_9740));
      --
    end process; 
    -- flow-through select operator MUX_9739_inst
    ISbox_in00_9740 <= IS00_9290 when (l_round_buffer(0) /=  '0') else IMX00_9599;
    -- logger for split-operator MUX_9745_inst flow-through 
    process(ISbox_in01_9746) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:MUX_9745_inst:flowthrough inputs: " & " l_round_buffer = "& Convert_SLV_To_Hex_String(l_round_buffer) & " IS01_9294 = "& Convert_SLV_To_Hex_String(IS01_9294) & " IMX01_9608 = "& Convert_SLV_To_Hex_String(IMX01_9608) & " outputs:" & " ISbox_in01_9746= "  & Convert_SLV_To_Hex_String(ISbox_in01_9746));
      --
    end process; 
    -- flow-through select operator MUX_9745_inst
    ISbox_in01_9746 <= IS01_9294 when (l_round_buffer(0) /=  '0') else IMX01_9608;
    -- logger for split-operator MUX_9751_inst flow-through 
    process(ISbox_in02_9752) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:MUX_9751_inst:flowthrough inputs: " & " l_round_buffer = "& Convert_SLV_To_Hex_String(l_round_buffer) & " IS02_9298 = "& Convert_SLV_To_Hex_String(IS02_9298) & " IMX02_9617 = "& Convert_SLV_To_Hex_String(IMX02_9617) & " outputs:" & " ISbox_in02_9752= "  & Convert_SLV_To_Hex_String(ISbox_in02_9752));
      --
    end process; 
    -- flow-through select operator MUX_9751_inst
    ISbox_in02_9752 <= IS02_9298 when (l_round_buffer(0) /=  '0') else IMX02_9617;
    -- logger for split-operator MUX_9757_inst flow-through 
    process(ISbox_in03_9758) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:MUX_9757_inst:flowthrough inputs: " & " l_round_buffer = "& Convert_SLV_To_Hex_String(l_round_buffer) & " IS03_9302 = "& Convert_SLV_To_Hex_String(IS03_9302) & " IMX03_9626 = "& Convert_SLV_To_Hex_String(IMX03_9626) & " outputs:" & " ISbox_in03_9758= "  & Convert_SLV_To_Hex_String(ISbox_in03_9758));
      --
    end process; 
    -- flow-through select operator MUX_9757_inst
    ISbox_in03_9758 <= IS03_9302 when (l_round_buffer(0) /=  '0') else IMX03_9626;
    -- logger for split-operator MUX_9763_inst flow-through 
    process(ISbox_in04_9764) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:MUX_9763_inst:flowthrough inputs: " & " l_round_buffer = "& Convert_SLV_To_Hex_String(l_round_buffer) & " IS04_9306 = "& Convert_SLV_To_Hex_String(IS04_9306) & " IMX04_9635 = "& Convert_SLV_To_Hex_String(IMX04_9635) & " outputs:" & " ISbox_in04_9764= "  & Convert_SLV_To_Hex_String(ISbox_in04_9764));
      --
    end process; 
    -- flow-through select operator MUX_9763_inst
    ISbox_in04_9764 <= IS04_9306 when (l_round_buffer(0) /=  '0') else IMX04_9635;
    -- logger for split-operator MUX_9769_inst flow-through 
    process(ISbox_in05_9770) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:MUX_9769_inst:flowthrough inputs: " & " l_round_buffer = "& Convert_SLV_To_Hex_String(l_round_buffer) & " IS05_9310 = "& Convert_SLV_To_Hex_String(IS05_9310) & " IMX05_9644 = "& Convert_SLV_To_Hex_String(IMX05_9644) & " outputs:" & " ISbox_in05_9770= "  & Convert_SLV_To_Hex_String(ISbox_in05_9770));
      --
    end process; 
    -- flow-through select operator MUX_9769_inst
    ISbox_in05_9770 <= IS05_9310 when (l_round_buffer(0) /=  '0') else IMX05_9644;
    -- logger for split-operator MUX_9775_inst flow-through 
    process(ISbox_in06_9776) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:MUX_9775_inst:flowthrough inputs: " & " l_round_buffer = "& Convert_SLV_To_Hex_String(l_round_buffer) & " IS06_9314 = "& Convert_SLV_To_Hex_String(IS06_9314) & " IMX06_9653 = "& Convert_SLV_To_Hex_String(IMX06_9653) & " outputs:" & " ISbox_in06_9776= "  & Convert_SLV_To_Hex_String(ISbox_in06_9776));
      --
    end process; 
    -- flow-through select operator MUX_9775_inst
    ISbox_in06_9776 <= IS06_9314 when (l_round_buffer(0) /=  '0') else IMX06_9653;
    -- logger for split-operator MUX_9781_inst flow-through 
    process(ISbox_in07_9782) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:MUX_9781_inst:flowthrough inputs: " & " l_round_buffer = "& Convert_SLV_To_Hex_String(l_round_buffer) & " IS07_9318 = "& Convert_SLV_To_Hex_String(IS07_9318) & " IMX07_9662 = "& Convert_SLV_To_Hex_String(IMX07_9662) & " outputs:" & " ISbox_in07_9782= "  & Convert_SLV_To_Hex_String(ISbox_in07_9782));
      --
    end process; 
    -- flow-through select operator MUX_9781_inst
    ISbox_in07_9782 <= IS07_9318 when (l_round_buffer(0) /=  '0') else IMX07_9662;
    -- logger for split-operator MUX_9787_inst flow-through 
    process(ISbox_in08_9788) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:MUX_9787_inst:flowthrough inputs: " & " l_round_buffer = "& Convert_SLV_To_Hex_String(l_round_buffer) & " IS08_9322 = "& Convert_SLV_To_Hex_String(IS08_9322) & " IMX08_9671 = "& Convert_SLV_To_Hex_String(IMX08_9671) & " outputs:" & " ISbox_in08_9788= "  & Convert_SLV_To_Hex_String(ISbox_in08_9788));
      --
    end process; 
    -- flow-through select operator MUX_9787_inst
    ISbox_in08_9788 <= IS08_9322 when (l_round_buffer(0) /=  '0') else IMX08_9671;
    -- logger for split-operator MUX_9793_inst flow-through 
    process(ISbox_in09_9794) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:MUX_9793_inst:flowthrough inputs: " & " l_round_buffer = "& Convert_SLV_To_Hex_String(l_round_buffer) & " IS09_9326 = "& Convert_SLV_To_Hex_String(IS09_9326) & " IMX09_9680 = "& Convert_SLV_To_Hex_String(IMX09_9680) & " outputs:" & " ISbox_in09_9794= "  & Convert_SLV_To_Hex_String(ISbox_in09_9794));
      --
    end process; 
    -- flow-through select operator MUX_9793_inst
    ISbox_in09_9794 <= IS09_9326 when (l_round_buffer(0) /=  '0') else IMX09_9680;
    -- logger for split-operator MUX_9799_inst flow-through 
    process(ISbox_in10_9800) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:MUX_9799_inst:flowthrough inputs: " & " l_round_buffer = "& Convert_SLV_To_Hex_String(l_round_buffer) & " IS10_9330 = "& Convert_SLV_To_Hex_String(IS10_9330) & " IMX10_9689 = "& Convert_SLV_To_Hex_String(IMX10_9689) & " outputs:" & " ISbox_in10_9800= "  & Convert_SLV_To_Hex_String(ISbox_in10_9800));
      --
    end process; 
    -- flow-through select operator MUX_9799_inst
    ISbox_in10_9800 <= IS10_9330 when (l_round_buffer(0) /=  '0') else IMX10_9689;
    -- logger for split-operator MUX_9805_inst flow-through 
    process(ISbox_in11_9806) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:MUX_9805_inst:flowthrough inputs: " & " l_round_buffer = "& Convert_SLV_To_Hex_String(l_round_buffer) & " IS11_9334 = "& Convert_SLV_To_Hex_String(IS11_9334) & " IMX11_9698 = "& Convert_SLV_To_Hex_String(IMX11_9698) & " outputs:" & " ISbox_in11_9806= "  & Convert_SLV_To_Hex_String(ISbox_in11_9806));
      --
    end process; 
    -- flow-through select operator MUX_9805_inst
    ISbox_in11_9806 <= IS11_9334 when (l_round_buffer(0) /=  '0') else IMX11_9698;
    -- logger for split-operator MUX_9811_inst flow-through 
    process(ISbox_in12_9812) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:MUX_9811_inst:flowthrough inputs: " & " l_round_buffer = "& Convert_SLV_To_Hex_String(l_round_buffer) & " IS12_9338 = "& Convert_SLV_To_Hex_String(IS12_9338) & " IMX12_9707 = "& Convert_SLV_To_Hex_String(IMX12_9707) & " outputs:" & " ISbox_in12_9812= "  & Convert_SLV_To_Hex_String(ISbox_in12_9812));
      --
    end process; 
    -- flow-through select operator MUX_9811_inst
    ISbox_in12_9812 <= IS12_9338 when (l_round_buffer(0) /=  '0') else IMX12_9707;
    -- logger for split-operator MUX_9817_inst flow-through 
    process(ISbox_in13_9818) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:MUX_9817_inst:flowthrough inputs: " & " l_round_buffer = "& Convert_SLV_To_Hex_String(l_round_buffer) & " IS13_9342 = "& Convert_SLV_To_Hex_String(IS13_9342) & " IMX13_9716 = "& Convert_SLV_To_Hex_String(IMX13_9716) & " outputs:" & " ISbox_in13_9818= "  & Convert_SLV_To_Hex_String(ISbox_in13_9818));
      --
    end process; 
    -- flow-through select operator MUX_9817_inst
    ISbox_in13_9818 <= IS13_9342 when (l_round_buffer(0) /=  '0') else IMX13_9716;
    -- logger for split-operator MUX_9823_inst flow-through 
    process(ISbox_in14_9824) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:MUX_9823_inst:flowthrough inputs: " & " l_round_buffer = "& Convert_SLV_To_Hex_String(l_round_buffer) & " IS14_9346 = "& Convert_SLV_To_Hex_String(IS14_9346) & " IMX14_9725 = "& Convert_SLV_To_Hex_String(IMX14_9725) & " outputs:" & " ISbox_in14_9824= "  & Convert_SLV_To_Hex_String(ISbox_in14_9824));
      --
    end process; 
    -- flow-through select operator MUX_9823_inst
    ISbox_in14_9824 <= IS14_9346 when (l_round_buffer(0) /=  '0') else IMX14_9725;
    -- logger for split-operator MUX_9829_inst flow-through 
    process(ISbox_in15_9830) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:MUX_9829_inst:flowthrough inputs: " & " l_round_buffer = "& Convert_SLV_To_Hex_String(l_round_buffer) & " IS15_9350 = "& Convert_SLV_To_Hex_String(IS15_9350) & " IMX15_9734 = "& Convert_SLV_To_Hex_String(IMX15_9734) & " outputs:" & " ISbox_in15_9830= "  & Convert_SLV_To_Hex_String(ISbox_in15_9830));
      --
    end process; 
    -- flow-through select operator MUX_9829_inst
    ISbox_in15_9830 <= IS15_9350 when (l_round_buffer(0) /=  '0') else IMX15_9734;
    -- logger for split-operator slice_9273_inst flow-through 
    process(ISa_9274) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:slice_9273_inst:flowthrough inputs: " & " round_in_buffer = "& Convert_SLV_To_Hex_String(round_in_buffer) & " outputs:" & " ISa_9274= "  & Convert_SLV_To_Hex_String(ISa_9274));
      --
    end process; 
    -- flow-through slice operator slice_9273_inst
    ISa_9274 <= round_in_buffer(127 downto 96);
    -- logger for split-operator slice_9277_inst flow-through 
    process(ISb_9278) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:slice_9277_inst:flowthrough inputs: " & " round_in_buffer = "& Convert_SLV_To_Hex_String(round_in_buffer) & " outputs:" & " ISb_9278= "  & Convert_SLV_To_Hex_String(ISb_9278));
      --
    end process; 
    -- flow-through slice operator slice_9277_inst
    ISb_9278 <= round_in_buffer(95 downto 64);
    -- logger for split-operator slice_9281_inst flow-through 
    process(ISc_9282) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:slice_9281_inst:flowthrough inputs: " & " round_in_buffer = "& Convert_SLV_To_Hex_String(round_in_buffer) & " outputs:" & " ISc_9282= "  & Convert_SLV_To_Hex_String(ISc_9282));
      --
    end process; 
    -- flow-through slice operator slice_9281_inst
    ISc_9282 <= round_in_buffer(63 downto 32);
    -- logger for split-operator slice_9285_inst flow-through 
    process(ISd_9286) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:slice_9285_inst:flowthrough inputs: " & " round_in_buffer = "& Convert_SLV_To_Hex_String(round_in_buffer) & " outputs:" & " ISd_9286= "  & Convert_SLV_To_Hex_String(ISd_9286));
      --
    end process; 
    -- flow-through slice operator slice_9285_inst
    ISd_9286 <= round_in_buffer(31 downto 0);
    -- logger for split-operator slice_9289_inst flow-through 
    process(IS00_9290) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:slice_9289_inst:flowthrough inputs: " & " ISa_9274 = "& Convert_SLV_To_Hex_String(ISa_9274) & " outputs:" & " IS00_9290= "  & Convert_SLV_To_Hex_String(IS00_9290));
      --
    end process; 
    -- flow-through slice operator slice_9289_inst
    IS00_9290 <= ISa_9274(31 downto 24);
    -- logger for split-operator slice_9293_inst flow-through 
    process(IS01_9294) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:slice_9293_inst:flowthrough inputs: " & " ISa_9274 = "& Convert_SLV_To_Hex_String(ISa_9274) & " outputs:" & " IS01_9294= "  & Convert_SLV_To_Hex_String(IS01_9294));
      --
    end process; 
    -- flow-through slice operator slice_9293_inst
    IS01_9294 <= ISa_9274(23 downto 16);
    -- logger for split-operator slice_9297_inst flow-through 
    process(IS02_9298) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:slice_9297_inst:flowthrough inputs: " & " ISa_9274 = "& Convert_SLV_To_Hex_String(ISa_9274) & " outputs:" & " IS02_9298= "  & Convert_SLV_To_Hex_String(IS02_9298));
      --
    end process; 
    -- flow-through slice operator slice_9297_inst
    IS02_9298 <= ISa_9274(15 downto 8);
    -- logger for split-operator slice_9301_inst flow-through 
    process(IS03_9302) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:slice_9301_inst:flowthrough inputs: " & " ISa_9274 = "& Convert_SLV_To_Hex_String(ISa_9274) & " outputs:" & " IS03_9302= "  & Convert_SLV_To_Hex_String(IS03_9302));
      --
    end process; 
    -- flow-through slice operator slice_9301_inst
    IS03_9302 <= ISa_9274(7 downto 0);
    -- logger for split-operator slice_9305_inst flow-through 
    process(IS04_9306) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:slice_9305_inst:flowthrough inputs: " & " ISb_9278 = "& Convert_SLV_To_Hex_String(ISb_9278) & " outputs:" & " IS04_9306= "  & Convert_SLV_To_Hex_String(IS04_9306));
      --
    end process; 
    -- flow-through slice operator slice_9305_inst
    IS04_9306 <= ISb_9278(31 downto 24);
    -- logger for split-operator slice_9309_inst flow-through 
    process(IS05_9310) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:slice_9309_inst:flowthrough inputs: " & " ISb_9278 = "& Convert_SLV_To_Hex_String(ISb_9278) & " outputs:" & " IS05_9310= "  & Convert_SLV_To_Hex_String(IS05_9310));
      --
    end process; 
    -- flow-through slice operator slice_9309_inst
    IS05_9310 <= ISb_9278(23 downto 16);
    -- logger for split-operator slice_9313_inst flow-through 
    process(IS06_9314) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:slice_9313_inst:flowthrough inputs: " & " ISb_9278 = "& Convert_SLV_To_Hex_String(ISb_9278) & " outputs:" & " IS06_9314= "  & Convert_SLV_To_Hex_String(IS06_9314));
      --
    end process; 
    -- flow-through slice operator slice_9313_inst
    IS06_9314 <= ISb_9278(15 downto 8);
    -- logger for split-operator slice_9317_inst flow-through 
    process(IS07_9318) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:slice_9317_inst:flowthrough inputs: " & " ISb_9278 = "& Convert_SLV_To_Hex_String(ISb_9278) & " outputs:" & " IS07_9318= "  & Convert_SLV_To_Hex_String(IS07_9318));
      --
    end process; 
    -- flow-through slice operator slice_9317_inst
    IS07_9318 <= ISb_9278(7 downto 0);
    -- logger for split-operator slice_9321_inst flow-through 
    process(IS08_9322) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:slice_9321_inst:flowthrough inputs: " & " ISc_9282 = "& Convert_SLV_To_Hex_String(ISc_9282) & " outputs:" & " IS08_9322= "  & Convert_SLV_To_Hex_String(IS08_9322));
      --
    end process; 
    -- flow-through slice operator slice_9321_inst
    IS08_9322 <= ISc_9282(31 downto 24);
    -- logger for split-operator slice_9325_inst flow-through 
    process(IS09_9326) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:slice_9325_inst:flowthrough inputs: " & " ISc_9282 = "& Convert_SLV_To_Hex_String(ISc_9282) & " outputs:" & " IS09_9326= "  & Convert_SLV_To_Hex_String(IS09_9326));
      --
    end process; 
    -- flow-through slice operator slice_9325_inst
    IS09_9326 <= ISc_9282(23 downto 16);
    -- logger for split-operator slice_9329_inst flow-through 
    process(IS10_9330) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:slice_9329_inst:flowthrough inputs: " & " ISc_9282 = "& Convert_SLV_To_Hex_String(ISc_9282) & " outputs:" & " IS10_9330= "  & Convert_SLV_To_Hex_String(IS10_9330));
      --
    end process; 
    -- flow-through slice operator slice_9329_inst
    IS10_9330 <= ISc_9282(15 downto 8);
    -- logger for split-operator slice_9333_inst flow-through 
    process(IS11_9334) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:slice_9333_inst:flowthrough inputs: " & " ISc_9282 = "& Convert_SLV_To_Hex_String(ISc_9282) & " outputs:" & " IS11_9334= "  & Convert_SLV_To_Hex_String(IS11_9334));
      --
    end process; 
    -- flow-through slice operator slice_9333_inst
    IS11_9334 <= ISc_9282(7 downto 0);
    -- logger for split-operator slice_9337_inst flow-through 
    process(IS12_9338) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:slice_9337_inst:flowthrough inputs: " & " ISd_9286 = "& Convert_SLV_To_Hex_String(ISd_9286) & " outputs:" & " IS12_9338= "  & Convert_SLV_To_Hex_String(IS12_9338));
      --
    end process; 
    -- flow-through slice operator slice_9337_inst
    IS12_9338 <= ISd_9286(31 downto 24);
    -- logger for split-operator slice_9341_inst flow-through 
    process(IS13_9342) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:slice_9341_inst:flowthrough inputs: " & " ISd_9286 = "& Convert_SLV_To_Hex_String(ISd_9286) & " outputs:" & " IS13_9342= "  & Convert_SLV_To_Hex_String(IS13_9342));
      --
    end process; 
    -- flow-through slice operator slice_9341_inst
    IS13_9342 <= ISd_9286(23 downto 16);
    -- logger for split-operator slice_9345_inst flow-through 
    process(IS14_9346) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:slice_9345_inst:flowthrough inputs: " & " ISd_9286 = "& Convert_SLV_To_Hex_String(ISd_9286) & " outputs:" & " IS14_9346= "  & Convert_SLV_To_Hex_String(IS14_9346));
      --
    end process; 
    -- flow-through slice operator slice_9345_inst
    IS14_9346 <= ISd_9286(15 downto 8);
    -- logger for split-operator slice_9349_inst flow-through 
    process(IS15_9350) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:slice_9349_inst:flowthrough inputs: " & " ISd_9286 = "& Convert_SLV_To_Hex_String(ISd_9286) & " outputs:" & " IS15_9350= "  & Convert_SLV_To_Hex_String(IS15_9350));
      --
    end process; 
    -- flow-through slice operator slice_9349_inst
    IS15_9350 <= ISd_9286(7 downto 0);
    -- logger for split-operator CONCAT_u16_u32_9886_inst flow-through 
    process(ISX0_9887) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:CONCAT_u16_u32_9886_inst:flowthrough inputs: " & " CONCAT_u8_u16_9882_wire = "& Convert_SLV_To_Hex_String(CONCAT_u8_u16_9882_wire) & " CONCAT_u8_u16_9885_wire = "& Convert_SLV_To_Hex_String(CONCAT_u8_u16_9885_wire) & " outputs:" & " ISX0_9887= "  & Convert_SLV_To_Hex_String(ISX0_9887));
      --
    end process; 
    -- binary operator CONCAT_u16_u32_9886_inst
    process(CONCAT_u8_u16_9882_wire, CONCAT_u8_u16_9885_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u8_u16_9882_wire, CONCAT_u8_u16_9885_wire, tmp_var);
      ISX0_9887 <= tmp_var; -- 
    end process;
    -- logger for split-operator CONCAT_u16_u32_9895_inst flow-through 
    process(ISX1_9896) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:CONCAT_u16_u32_9895_inst:flowthrough inputs: " & " CONCAT_u8_u16_9891_wire = "& Convert_SLV_To_Hex_String(CONCAT_u8_u16_9891_wire) & " CONCAT_u8_u16_9894_wire = "& Convert_SLV_To_Hex_String(CONCAT_u8_u16_9894_wire) & " outputs:" & " ISX1_9896= "  & Convert_SLV_To_Hex_String(ISX1_9896));
      --
    end process; 
    -- binary operator CONCAT_u16_u32_9895_inst
    process(CONCAT_u8_u16_9891_wire, CONCAT_u8_u16_9894_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u8_u16_9891_wire, CONCAT_u8_u16_9894_wire, tmp_var);
      ISX1_9896 <= tmp_var; -- 
    end process;
    -- logger for split-operator CONCAT_u16_u32_9904_inst flow-through 
    process(ISX2_9905) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:CONCAT_u16_u32_9904_inst:flowthrough inputs: " & " CONCAT_u8_u16_9900_wire = "& Convert_SLV_To_Hex_String(CONCAT_u8_u16_9900_wire) & " CONCAT_u8_u16_9903_wire = "& Convert_SLV_To_Hex_String(CONCAT_u8_u16_9903_wire) & " outputs:" & " ISX2_9905= "  & Convert_SLV_To_Hex_String(ISX2_9905));
      --
    end process; 
    -- binary operator CONCAT_u16_u32_9904_inst
    process(CONCAT_u8_u16_9900_wire, CONCAT_u8_u16_9903_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u8_u16_9900_wire, CONCAT_u8_u16_9903_wire, tmp_var);
      ISX2_9905 <= tmp_var; -- 
    end process;
    -- logger for split-operator CONCAT_u16_u32_9913_inst flow-through 
    process(ISX3_9914) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:CONCAT_u16_u32_9913_inst:flowthrough inputs: " & " CONCAT_u8_u16_9909_wire = "& Convert_SLV_To_Hex_String(CONCAT_u8_u16_9909_wire) & " CONCAT_u8_u16_9912_wire = "& Convert_SLV_To_Hex_String(CONCAT_u8_u16_9912_wire) & " outputs:" & " ISX3_9914= "  & Convert_SLV_To_Hex_String(ISX3_9914));
      --
    end process; 
    -- binary operator CONCAT_u16_u32_9913_inst
    process(CONCAT_u8_u16_9909_wire, CONCAT_u8_u16_9912_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u8_u16_9909_wire, CONCAT_u8_u16_9912_wire, tmp_var);
      ISX3_9914 <= tmp_var; -- 
    end process;
    -- logger for split-operator CONCAT_u32_u64_9918_inst flow-through 
    process(CONCAT_u32_u64_9918_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:CONCAT_u32_u64_9918_inst:flowthrough inputs: " & " ISX0_9887 = "& Convert_SLV_To_Hex_String(ISX0_9887) & " ISX1_9896 = "& Convert_SLV_To_Hex_String(ISX1_9896) & " outputs:" & " CONCAT_u32_u64_9918_wire= "  & Convert_SLV_To_Hex_String(CONCAT_u32_u64_9918_wire));
      --
    end process; 
    -- binary operator CONCAT_u32_u64_9918_inst
    process(ISX0_9887, ISX1_9896) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApConcat_proc(ISX0_9887, ISX1_9896, tmp_var);
      CONCAT_u32_u64_9918_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator CONCAT_u32_u64_9921_inst flow-through 
    process(CONCAT_u32_u64_9921_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:CONCAT_u32_u64_9921_inst:flowthrough inputs: " & " ISX2_9905 = "& Convert_SLV_To_Hex_String(ISX2_9905) & " ISX3_9914 = "& Convert_SLV_To_Hex_String(ISX3_9914) & " outputs:" & " CONCAT_u32_u64_9921_wire= "  & Convert_SLV_To_Hex_String(CONCAT_u32_u64_9921_wire));
      --
    end process; 
    -- binary operator CONCAT_u32_u64_9921_inst
    process(ISX2_9905, ISX3_9914) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApConcat_proc(ISX2_9905, ISX3_9914, tmp_var);
      CONCAT_u32_u64_9921_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator CONCAT_u64_u128_9922_inst flow-through 
    process(OUT_9923) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:CONCAT_u64_u128_9922_inst:flowthrough inputs: " & " CONCAT_u32_u64_9918_wire = "& Convert_SLV_To_Hex_String(CONCAT_u32_u64_9918_wire) & " CONCAT_u32_u64_9921_wire = "& Convert_SLV_To_Hex_String(CONCAT_u32_u64_9921_wire) & " outputs:" & " OUT_9923= "  & Convert_SLV_To_Hex_String(OUT_9923));
      --
    end process; 
    -- binary operator CONCAT_u64_u128_9922_inst
    process(CONCAT_u32_u64_9918_wire, CONCAT_u32_u64_9921_wire) -- 
      variable tmp_var : std_logic_vector(127 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u32_u64_9918_wire, CONCAT_u32_u64_9921_wire, tmp_var);
      OUT_9923 <= tmp_var; -- 
    end process;
    -- logger for split-operator CONCAT_u8_u16_9882_inst flow-through 
    process(CONCAT_u8_u16_9882_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:CONCAT_u8_u16_9882_inst:flowthrough inputs: " & " Sout00_9833 = "& Convert_SLV_To_Hex_String(Sout00_9833) & " Sout01_9872 = "& Convert_SLV_To_Hex_String(Sout01_9872) & " outputs:" & " CONCAT_u8_u16_9882_wire= "  & Convert_SLV_To_Hex_String(CONCAT_u8_u16_9882_wire));
      --
    end process; 
    -- binary operator CONCAT_u8_u16_9882_inst
    process(Sout00_9833, Sout01_9872) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApConcat_proc(Sout00_9833, Sout01_9872, tmp_var);
      CONCAT_u8_u16_9882_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator CONCAT_u8_u16_9885_inst flow-through 
    process(CONCAT_u8_u16_9885_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:CONCAT_u8_u16_9885_inst:flowthrough inputs: " & " Sout02_9863 = "& Convert_SLV_To_Hex_String(Sout02_9863) & " Sout03_9854 = "& Convert_SLV_To_Hex_String(Sout03_9854) & " outputs:" & " CONCAT_u8_u16_9885_wire= "  & Convert_SLV_To_Hex_String(CONCAT_u8_u16_9885_wire));
      --
    end process; 
    -- binary operator CONCAT_u8_u16_9885_inst
    process(Sout02_9863, Sout03_9854) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApConcat_proc(Sout02_9863, Sout03_9854, tmp_var);
      CONCAT_u8_u16_9885_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator CONCAT_u8_u16_9891_inst flow-through 
    process(CONCAT_u8_u16_9891_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:CONCAT_u8_u16_9891_inst:flowthrough inputs: " & " Sout04_9845 = "& Convert_SLV_To_Hex_String(Sout04_9845) & " Sout05_9836 = "& Convert_SLV_To_Hex_String(Sout05_9836) & " outputs:" & " CONCAT_u8_u16_9891_wire= "  & Convert_SLV_To_Hex_String(CONCAT_u8_u16_9891_wire));
      --
    end process; 
    -- binary operator CONCAT_u8_u16_9891_inst
    process(Sout04_9845, Sout05_9836) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApConcat_proc(Sout04_9845, Sout05_9836, tmp_var);
      CONCAT_u8_u16_9891_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator CONCAT_u8_u16_9894_inst flow-through 
    process(CONCAT_u8_u16_9894_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:CONCAT_u8_u16_9894_inst:flowthrough inputs: " & " Sout06_9875 = "& Convert_SLV_To_Hex_String(Sout06_9875) & " Sout07_9866 = "& Convert_SLV_To_Hex_String(Sout07_9866) & " outputs:" & " CONCAT_u8_u16_9894_wire= "  & Convert_SLV_To_Hex_String(CONCAT_u8_u16_9894_wire));
      --
    end process; 
    -- binary operator CONCAT_u8_u16_9894_inst
    process(Sout06_9875, Sout07_9866) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApConcat_proc(Sout06_9875, Sout07_9866, tmp_var);
      CONCAT_u8_u16_9894_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator CONCAT_u8_u16_9900_inst flow-through 
    process(CONCAT_u8_u16_9900_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:CONCAT_u8_u16_9900_inst:flowthrough inputs: " & " Sout08_9857 = "& Convert_SLV_To_Hex_String(Sout08_9857) & " Sout09_9848 = "& Convert_SLV_To_Hex_String(Sout09_9848) & " outputs:" & " CONCAT_u8_u16_9900_wire= "  & Convert_SLV_To_Hex_String(CONCAT_u8_u16_9900_wire));
      --
    end process; 
    -- binary operator CONCAT_u8_u16_9900_inst
    process(Sout08_9857, Sout09_9848) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApConcat_proc(Sout08_9857, Sout09_9848, tmp_var);
      CONCAT_u8_u16_9900_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator CONCAT_u8_u16_9903_inst flow-through 
    process(CONCAT_u8_u16_9903_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:CONCAT_u8_u16_9903_inst:flowthrough inputs: " & " Sout10_9839 = "& Convert_SLV_To_Hex_String(Sout10_9839) & " Sout11_9878 = "& Convert_SLV_To_Hex_String(Sout11_9878) & " outputs:" & " CONCAT_u8_u16_9903_wire= "  & Convert_SLV_To_Hex_String(CONCAT_u8_u16_9903_wire));
      --
    end process; 
    -- binary operator CONCAT_u8_u16_9903_inst
    process(Sout10_9839, Sout11_9878) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApConcat_proc(Sout10_9839, Sout11_9878, tmp_var);
      CONCAT_u8_u16_9903_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator CONCAT_u8_u16_9909_inst flow-through 
    process(CONCAT_u8_u16_9909_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:CONCAT_u8_u16_9909_inst:flowthrough inputs: " & " Sout12_9869 = "& Convert_SLV_To_Hex_String(Sout12_9869) & " Sout13_9860 = "& Convert_SLV_To_Hex_String(Sout13_9860) & " outputs:" & " CONCAT_u8_u16_9909_wire= "  & Convert_SLV_To_Hex_String(CONCAT_u8_u16_9909_wire));
      --
    end process; 
    -- binary operator CONCAT_u8_u16_9909_inst
    process(Sout12_9869, Sout13_9860) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApConcat_proc(Sout12_9869, Sout13_9860, tmp_var);
      CONCAT_u8_u16_9909_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator CONCAT_u8_u16_9912_inst flow-through 
    process(CONCAT_u8_u16_9912_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:CONCAT_u8_u16_9912_inst:flowthrough inputs: " & " Sout14_9851 = "& Convert_SLV_To_Hex_String(Sout14_9851) & " Sout15_9842 = "& Convert_SLV_To_Hex_String(Sout15_9842) & " outputs:" & " CONCAT_u8_u16_9912_wire= "  & Convert_SLV_To_Hex_String(CONCAT_u8_u16_9912_wire));
      --
    end process; 
    -- binary operator CONCAT_u8_u16_9912_inst
    process(Sout14_9851, Sout15_9842) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApConcat_proc(Sout14_9851, Sout15_9842, tmp_var);
      CONCAT_u8_u16_9912_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator XOR_u128_u128_9927_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if XOR_u128_u128_9927_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:XOR_u128_u128_9927_inst:started:   inputs: " & " OUT_9923 = "& Convert_SLV_To_Hex_String(OUT_9923) & " key_in_buffer = "& Convert_SLV_To_Hex_String(key_in_buffer));
          --
        end if; 
        if XOR_u128_u128_9927_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:XOR_u128_u128_9927_inst:finished:  outputs: " & " round_out_buffer= "  & Convert_SLV_To_Hex_String(round_out_buffer));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (15) : XOR_u128_u128_9927_inst 
    ApIntXor_group_15: Block -- 
      signal data_in: std_logic_vector(255 downto 0);
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= OUT_9923 & key_in_buffer;
      round_out_buffer <= data_out(127 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= XOR_u128_u128_9927_inst_req_0;
      XOR_u128_u128_9927_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= XOR_u128_u128_9927_inst_req_1;
      XOR_u128_u128_9927_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntXor",
          name => "ApIntXor_group_15",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 128,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 128, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 128,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 15
    -- logger for split-operator XOR_u8_u8_9402_inst flow-through 
    process(XOR_u8_u8_9402_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:XOR_u8_u8_9402_inst:flowthrough inputs: " & " IS00_9290 = "& Convert_SLV_To_Hex_String(IS00_9290) & " IS01_9294 = "& Convert_SLV_To_Hex_String(IS01_9294) & " outputs:" & " XOR_u8_u8_9402_wire= "  & Convert_SLV_To_Hex_String(XOR_u8_u8_9402_wire));
      --
    end process; 
    -- binary operator XOR_u8_u8_9402_inst
    process(IS00_9290, IS01_9294) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(IS00_9290, IS01_9294, tmp_var);
      XOR_u8_u8_9402_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator XOR_u8_u8_9405_inst flow-through 
    process(XOR_u8_u8_9405_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:XOR_u8_u8_9405_inst:flowthrough inputs: " & " IS02_9298 = "& Convert_SLV_To_Hex_String(IS02_9298) & " IS03_9302 = "& Convert_SLV_To_Hex_String(IS03_9302) & " outputs:" & " XOR_u8_u8_9405_wire= "  & Convert_SLV_To_Hex_String(XOR_u8_u8_9405_wire));
      --
    end process; 
    -- binary operator XOR_u8_u8_9405_inst
    process(IS02_9298, IS03_9302) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(IS02_9298, IS03_9302, tmp_var);
      XOR_u8_u8_9405_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator XOR_u8_u8_9406_inst flow-through 
    process(Wc0_9407) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:XOR_u8_u8_9406_inst:flowthrough inputs: " & " XOR_u8_u8_9402_wire = "& Convert_SLV_To_Hex_String(XOR_u8_u8_9402_wire) & " XOR_u8_u8_9405_wire = "& Convert_SLV_To_Hex_String(XOR_u8_u8_9405_wire) & " outputs:" & " Wc0_9407= "  & Convert_SLV_To_Hex_String(Wc0_9407));
      --
    end process; 
    -- binary operator XOR_u8_u8_9406_inst
    process(XOR_u8_u8_9402_wire, XOR_u8_u8_9405_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(XOR_u8_u8_9402_wire, XOR_u8_u8_9405_wire, tmp_var);
      Wc0_9407 <= tmp_var; -- 
    end process;
    -- logger for split-operator XOR_u8_u8_9411_inst flow-through 
    process(XOR_u8_u8_9411_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:XOR_u8_u8_9411_inst:flowthrough inputs: " & " IS04_9306 = "& Convert_SLV_To_Hex_String(IS04_9306) & " IS05_9310 = "& Convert_SLV_To_Hex_String(IS05_9310) & " outputs:" & " XOR_u8_u8_9411_wire= "  & Convert_SLV_To_Hex_String(XOR_u8_u8_9411_wire));
      --
    end process; 
    -- binary operator XOR_u8_u8_9411_inst
    process(IS04_9306, IS05_9310) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(IS04_9306, IS05_9310, tmp_var);
      XOR_u8_u8_9411_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator XOR_u8_u8_9414_inst flow-through 
    process(XOR_u8_u8_9414_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:XOR_u8_u8_9414_inst:flowthrough inputs: " & " IS06_9314 = "& Convert_SLV_To_Hex_String(IS06_9314) & " IS07_9318 = "& Convert_SLV_To_Hex_String(IS07_9318) & " outputs:" & " XOR_u8_u8_9414_wire= "  & Convert_SLV_To_Hex_String(XOR_u8_u8_9414_wire));
      --
    end process; 
    -- binary operator XOR_u8_u8_9414_inst
    process(IS06_9314, IS07_9318) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(IS06_9314, IS07_9318, tmp_var);
      XOR_u8_u8_9414_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator XOR_u8_u8_9415_inst flow-through 
    process(Wc1_9416) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:XOR_u8_u8_9415_inst:flowthrough inputs: " & " XOR_u8_u8_9411_wire = "& Convert_SLV_To_Hex_String(XOR_u8_u8_9411_wire) & " XOR_u8_u8_9414_wire = "& Convert_SLV_To_Hex_String(XOR_u8_u8_9414_wire) & " outputs:" & " Wc1_9416= "  & Convert_SLV_To_Hex_String(Wc1_9416));
      --
    end process; 
    -- binary operator XOR_u8_u8_9415_inst
    process(XOR_u8_u8_9411_wire, XOR_u8_u8_9414_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(XOR_u8_u8_9411_wire, XOR_u8_u8_9414_wire, tmp_var);
      Wc1_9416 <= tmp_var; -- 
    end process;
    -- logger for split-operator XOR_u8_u8_9420_inst flow-through 
    process(XOR_u8_u8_9420_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:XOR_u8_u8_9420_inst:flowthrough inputs: " & " IS08_9322 = "& Convert_SLV_To_Hex_String(IS08_9322) & " IS09_9326 = "& Convert_SLV_To_Hex_String(IS09_9326) & " outputs:" & " XOR_u8_u8_9420_wire= "  & Convert_SLV_To_Hex_String(XOR_u8_u8_9420_wire));
      --
    end process; 
    -- binary operator XOR_u8_u8_9420_inst
    process(IS08_9322, IS09_9326) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(IS08_9322, IS09_9326, tmp_var);
      XOR_u8_u8_9420_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator XOR_u8_u8_9423_inst flow-through 
    process(XOR_u8_u8_9423_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:XOR_u8_u8_9423_inst:flowthrough inputs: " & " IS10_9330 = "& Convert_SLV_To_Hex_String(IS10_9330) & " IS11_9334 = "& Convert_SLV_To_Hex_String(IS11_9334) & " outputs:" & " XOR_u8_u8_9423_wire= "  & Convert_SLV_To_Hex_String(XOR_u8_u8_9423_wire));
      --
    end process; 
    -- binary operator XOR_u8_u8_9423_inst
    process(IS10_9330, IS11_9334) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(IS10_9330, IS11_9334, tmp_var);
      XOR_u8_u8_9423_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator XOR_u8_u8_9424_inst flow-through 
    process(Wc2_9425) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:XOR_u8_u8_9424_inst:flowthrough inputs: " & " XOR_u8_u8_9420_wire = "& Convert_SLV_To_Hex_String(XOR_u8_u8_9420_wire) & " XOR_u8_u8_9423_wire = "& Convert_SLV_To_Hex_String(XOR_u8_u8_9423_wire) & " outputs:" & " Wc2_9425= "  & Convert_SLV_To_Hex_String(Wc2_9425));
      --
    end process; 
    -- binary operator XOR_u8_u8_9424_inst
    process(XOR_u8_u8_9420_wire, XOR_u8_u8_9423_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(XOR_u8_u8_9420_wire, XOR_u8_u8_9423_wire, tmp_var);
      Wc2_9425 <= tmp_var; -- 
    end process;
    -- logger for split-operator XOR_u8_u8_9429_inst flow-through 
    process(XOR_u8_u8_9429_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:XOR_u8_u8_9429_inst:flowthrough inputs: " & " IS12_9338 = "& Convert_SLV_To_Hex_String(IS12_9338) & " IS13_9342 = "& Convert_SLV_To_Hex_String(IS13_9342) & " outputs:" & " XOR_u8_u8_9429_wire= "  & Convert_SLV_To_Hex_String(XOR_u8_u8_9429_wire));
      --
    end process; 
    -- binary operator XOR_u8_u8_9429_inst
    process(IS12_9338, IS13_9342) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(IS12_9338, IS13_9342, tmp_var);
      XOR_u8_u8_9429_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator XOR_u8_u8_9432_inst flow-through 
    process(XOR_u8_u8_9432_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:XOR_u8_u8_9432_inst:flowthrough inputs: " & " IS14_9346 = "& Convert_SLV_To_Hex_String(IS14_9346) & " IS15_9350 = "& Convert_SLV_To_Hex_String(IS15_9350) & " outputs:" & " XOR_u8_u8_9432_wire= "  & Convert_SLV_To_Hex_String(XOR_u8_u8_9432_wire));
      --
    end process; 
    -- binary operator XOR_u8_u8_9432_inst
    process(IS14_9346, IS15_9350) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(IS14_9346, IS15_9350, tmp_var);
      XOR_u8_u8_9432_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator XOR_u8_u8_9433_inst flow-through 
    process(Wc3_9434) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:XOR_u8_u8_9433_inst:flowthrough inputs: " & " XOR_u8_u8_9429_wire = "& Convert_SLV_To_Hex_String(XOR_u8_u8_9429_wire) & " XOR_u8_u8_9432_wire = "& Convert_SLV_To_Hex_String(XOR_u8_u8_9432_wire) & " outputs:" & " Wc3_9434= "  & Convert_SLV_To_Hex_String(Wc3_9434));
      --
    end process; 
    -- binary operator XOR_u8_u8_9433_inst
    process(XOR_u8_u8_9429_wire, XOR_u8_u8_9432_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(XOR_u8_u8_9429_wire, XOR_u8_u8_9432_wire, tmp_var);
      Wc3_9434 <= tmp_var; -- 
    end process;
    -- logger for split-operator XOR_u8_u8_9438_inst flow-through 
    process(Y00_9439) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:XOR_u8_u8_9438_inst:flowthrough inputs: " & " IS00x2_9353 = "& Convert_SLV_To_Hex_String(IS00x2_9353) & " IS02x2_9359 = "& Convert_SLV_To_Hex_String(IS02x2_9359) & " outputs:" & " Y00_9439= "  & Convert_SLV_To_Hex_String(Y00_9439));
      --
    end process; 
    -- binary operator XOR_u8_u8_9438_inst
    process(IS00x2_9353, IS02x2_9359) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(IS00x2_9353, IS02x2_9359, tmp_var);
      Y00_9439 <= tmp_var; -- 
    end process;
    -- logger for split-operator XOR_u8_u8_9443_inst flow-through 
    process(Y01_9444) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:XOR_u8_u8_9443_inst:flowthrough inputs: " & " IS04x2_9365 = "& Convert_SLV_To_Hex_String(IS04x2_9365) & " IS06x2_9371 = "& Convert_SLV_To_Hex_String(IS06x2_9371) & " outputs:" & " Y01_9444= "  & Convert_SLV_To_Hex_String(Y01_9444));
      --
    end process; 
    -- binary operator XOR_u8_u8_9443_inst
    process(IS04x2_9365, IS06x2_9371) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(IS04x2_9365, IS06x2_9371, tmp_var);
      Y01_9444 <= tmp_var; -- 
    end process;
    -- logger for split-operator XOR_u8_u8_9448_inst flow-through 
    process(Y02_9449) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:XOR_u8_u8_9448_inst:flowthrough inputs: " & " IS08x2_9377 = "& Convert_SLV_To_Hex_String(IS08x2_9377) & " IS10x2_9383 = "& Convert_SLV_To_Hex_String(IS10x2_9383) & " outputs:" & " Y02_9449= "  & Convert_SLV_To_Hex_String(Y02_9449));
      --
    end process; 
    -- binary operator XOR_u8_u8_9448_inst
    process(IS08x2_9377, IS10x2_9383) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(IS08x2_9377, IS10x2_9383, tmp_var);
      Y02_9449 <= tmp_var; -- 
    end process;
    -- logger for split-operator XOR_u8_u8_9453_inst flow-through 
    process(Y03_9454) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:XOR_u8_u8_9453_inst:flowthrough inputs: " & " IS12x2_9389 = "& Convert_SLV_To_Hex_String(IS12x2_9389) & " IS14x2_9395 = "& Convert_SLV_To_Hex_String(IS14x2_9395) & " outputs:" & " Y03_9454= "  & Convert_SLV_To_Hex_String(Y03_9454));
      --
    end process; 
    -- binary operator XOR_u8_u8_9453_inst
    process(IS12x2_9389, IS14x2_9395) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(IS12x2_9389, IS14x2_9395, tmp_var);
      Y03_9454 <= tmp_var; -- 
    end process;
    -- logger for split-operator XOR_u8_u8_9458_inst flow-through 
    process(Y10_9459) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:XOR_u8_u8_9458_inst:flowthrough inputs: " & " IS01x2_9356 = "& Convert_SLV_To_Hex_String(IS01x2_9356) & " IS03x2_9362 = "& Convert_SLV_To_Hex_String(IS03x2_9362) & " outputs:" & " Y10_9459= "  & Convert_SLV_To_Hex_String(Y10_9459));
      --
    end process; 
    -- binary operator XOR_u8_u8_9458_inst
    process(IS01x2_9356, IS03x2_9362) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(IS01x2_9356, IS03x2_9362, tmp_var);
      Y10_9459 <= tmp_var; -- 
    end process;
    -- logger for split-operator XOR_u8_u8_9463_inst flow-through 
    process(Y11_9464) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:XOR_u8_u8_9463_inst:flowthrough inputs: " & " IS05x2_9368 = "& Convert_SLV_To_Hex_String(IS05x2_9368) & " IS07x2_9374 = "& Convert_SLV_To_Hex_String(IS07x2_9374) & " outputs:" & " Y11_9464= "  & Convert_SLV_To_Hex_String(Y11_9464));
      --
    end process; 
    -- binary operator XOR_u8_u8_9463_inst
    process(IS05x2_9368, IS07x2_9374) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(IS05x2_9368, IS07x2_9374, tmp_var);
      Y11_9464 <= tmp_var; -- 
    end process;
    -- logger for split-operator XOR_u8_u8_9468_inst flow-through 
    process(Y12_9469) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:XOR_u8_u8_9468_inst:flowthrough inputs: " & " IS09x2_9380 = "& Convert_SLV_To_Hex_String(IS09x2_9380) & " IS11x2_9386 = "& Convert_SLV_To_Hex_String(IS11x2_9386) & " outputs:" & " Y12_9469= "  & Convert_SLV_To_Hex_String(Y12_9469));
      --
    end process; 
    -- binary operator XOR_u8_u8_9468_inst
    process(IS09x2_9380, IS11x2_9386) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(IS09x2_9380, IS11x2_9386, tmp_var);
      Y12_9469 <= tmp_var; -- 
    end process;
    -- logger for split-operator XOR_u8_u8_9473_inst flow-through 
    process(Y13_9474) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:XOR_u8_u8_9473_inst:flowthrough inputs: " & " IS13x2_9392 = "& Convert_SLV_To_Hex_String(IS13x2_9392) & " IS15x2_9398 = "& Convert_SLV_To_Hex_String(IS15x2_9398) & " outputs:" & " Y13_9474= "  & Convert_SLV_To_Hex_String(Y13_9474));
      --
    end process; 
    -- binary operator XOR_u8_u8_9473_inst
    process(IS13x2_9392, IS15x2_9398) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(IS13x2_9392, IS15x2_9398, tmp_var);
      Y13_9474 <= tmp_var; -- 
    end process;
    -- logger for split-operator XOR_u8_u8_9502_inst flow-through 
    process(Z0_9503) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:XOR_u8_u8_9502_inst:flowthrough inputs: " & " Y00x2_9477 = "& Convert_SLV_To_Hex_String(Y00x2_9477) & " Y10x2_9489 = "& Convert_SLV_To_Hex_String(Y10x2_9489) & " outputs:" & " Z0_9503= "  & Convert_SLV_To_Hex_String(Z0_9503));
      --
    end process; 
    -- binary operator XOR_u8_u8_9502_inst
    process(Y00x2_9477, Y10x2_9489) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(Y00x2_9477, Y10x2_9489, tmp_var);
      Z0_9503 <= tmp_var; -- 
    end process;
    -- logger for split-operator XOR_u8_u8_9507_inst flow-through 
    process(Z1_9508) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:XOR_u8_u8_9507_inst:flowthrough inputs: " & " Y01x2_9480 = "& Convert_SLV_To_Hex_String(Y01x2_9480) & " Y11x2_9492 = "& Convert_SLV_To_Hex_String(Y11x2_9492) & " outputs:" & " Z1_9508= "  & Convert_SLV_To_Hex_String(Z1_9508));
      --
    end process; 
    -- binary operator XOR_u8_u8_9507_inst
    process(Y01x2_9480, Y11x2_9492) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(Y01x2_9480, Y11x2_9492, tmp_var);
      Z1_9508 <= tmp_var; -- 
    end process;
    -- logger for split-operator XOR_u8_u8_9512_inst flow-through 
    process(Z2_9513) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:XOR_u8_u8_9512_inst:flowthrough inputs: " & " Y02x2_9483 = "& Convert_SLV_To_Hex_String(Y02x2_9483) & " Y12x2_9495 = "& Convert_SLV_To_Hex_String(Y12x2_9495) & " outputs:" & " Z2_9513= "  & Convert_SLV_To_Hex_String(Z2_9513));
      --
    end process; 
    -- binary operator XOR_u8_u8_9512_inst
    process(Y02x2_9483, Y12x2_9495) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(Y02x2_9483, Y12x2_9495, tmp_var);
      Z2_9513 <= tmp_var; -- 
    end process;
    -- logger for split-operator XOR_u8_u8_9517_inst flow-through 
    process(Z3_9518) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:XOR_u8_u8_9517_inst:flowthrough inputs: " & " Y03x2_9486 = "& Convert_SLV_To_Hex_String(Y03x2_9486) & " Y13x2_9498 = "& Convert_SLV_To_Hex_String(Y13x2_9498) & " outputs:" & " Z3_9518= "  & Convert_SLV_To_Hex_String(Z3_9518));
      --
    end process; 
    -- binary operator XOR_u8_u8_9517_inst
    process(Y03x2_9486, Y13x2_9498) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(Y03x2_9486, Y13x2_9498, tmp_var);
      Z3_9518 <= tmp_var; -- 
    end process;
    -- logger for split-operator XOR_u8_u8_9534_inst flow-through 
    process(A0_9535) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:XOR_u8_u8_9534_inst:flowthrough inputs: " & " Z0x2_9521 = "& Convert_SLV_To_Hex_String(Z0x2_9521) & " Wc0_9407 = "& Convert_SLV_To_Hex_String(Wc0_9407) & " outputs:" & " A0_9535= "  & Convert_SLV_To_Hex_String(A0_9535));
      --
    end process; 
    -- binary operator XOR_u8_u8_9534_inst
    process(Z0x2_9521, Wc0_9407) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(Z0x2_9521, Wc0_9407, tmp_var);
      A0_9535 <= tmp_var; -- 
    end process;
    -- logger for split-operator XOR_u8_u8_9539_inst flow-through 
    process(A1_9540) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:XOR_u8_u8_9539_inst:flowthrough inputs: " & " Z1x2_9524 = "& Convert_SLV_To_Hex_String(Z1x2_9524) & " Wc1_9416 = "& Convert_SLV_To_Hex_String(Wc1_9416) & " outputs:" & " A1_9540= "  & Convert_SLV_To_Hex_String(A1_9540));
      --
    end process; 
    -- binary operator XOR_u8_u8_9539_inst
    process(Z1x2_9524, Wc1_9416) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(Z1x2_9524, Wc1_9416, tmp_var);
      A1_9540 <= tmp_var; -- 
    end process;
    -- logger for split-operator XOR_u8_u8_9544_inst flow-through 
    process(A2_9545) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:XOR_u8_u8_9544_inst:flowthrough inputs: " & " Z2x2_9527 = "& Convert_SLV_To_Hex_String(Z2x2_9527) & " Wc2_9425 = "& Convert_SLV_To_Hex_String(Wc2_9425) & " outputs:" & " A2_9545= "  & Convert_SLV_To_Hex_String(A2_9545));
      --
    end process; 
    -- binary operator XOR_u8_u8_9544_inst
    process(Z2x2_9527, Wc2_9425) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(Z2x2_9527, Wc2_9425, tmp_var);
      A2_9545 <= tmp_var; -- 
    end process;
    -- logger for split-operator XOR_u8_u8_9549_inst flow-through 
    process(A3_9550) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:XOR_u8_u8_9549_inst:flowthrough inputs: " & " Z3x2_9530 = "& Convert_SLV_To_Hex_String(Z3x2_9530) & " Wc3_9434 = "& Convert_SLV_To_Hex_String(Wc3_9434) & " outputs:" & " A3_9550= "  & Convert_SLV_To_Hex_String(A3_9550));
      --
    end process; 
    -- binary operator XOR_u8_u8_9549_inst
    process(Z3x2_9530, Wc3_9434) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(Z3x2_9530, Wc3_9434, tmp_var);
      A3_9550 <= tmp_var; -- 
    end process;
    -- logger for split-operator XOR_u8_u8_9554_inst flow-through 
    process(B00_9555) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:XOR_u8_u8_9554_inst:flowthrough inputs: " & " A0_9535 = "& Convert_SLV_To_Hex_String(A0_9535) & " Y00x2_9477 = "& Convert_SLV_To_Hex_String(Y00x2_9477) & " outputs:" & " B00_9555= "  & Convert_SLV_To_Hex_String(B00_9555));
      --
    end process; 
    -- binary operator XOR_u8_u8_9554_inst
    process(A0_9535, Y00x2_9477) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(A0_9535, Y00x2_9477, tmp_var);
      B00_9555 <= tmp_var; -- 
    end process;
    -- logger for split-operator XOR_u8_u8_9559_inst flow-through 
    process(B01_9560) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:XOR_u8_u8_9559_inst:flowthrough inputs: " & " A1_9540 = "& Convert_SLV_To_Hex_String(A1_9540) & " Y01x2_9480 = "& Convert_SLV_To_Hex_String(Y01x2_9480) & " outputs:" & " B01_9560= "  & Convert_SLV_To_Hex_String(B01_9560));
      --
    end process; 
    -- binary operator XOR_u8_u8_9559_inst
    process(A1_9540, Y01x2_9480) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(A1_9540, Y01x2_9480, tmp_var);
      B01_9560 <= tmp_var; -- 
    end process;
    -- logger for split-operator XOR_u8_u8_9564_inst flow-through 
    process(B02_9565) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:XOR_u8_u8_9564_inst:flowthrough inputs: " & " A2_9545 = "& Convert_SLV_To_Hex_String(A2_9545) & " Y02x2_9483 = "& Convert_SLV_To_Hex_String(Y02x2_9483) & " outputs:" & " B02_9565= "  & Convert_SLV_To_Hex_String(B02_9565));
      --
    end process; 
    -- binary operator XOR_u8_u8_9564_inst
    process(A2_9545, Y02x2_9483) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(A2_9545, Y02x2_9483, tmp_var);
      B02_9565 <= tmp_var; -- 
    end process;
    -- logger for split-operator XOR_u8_u8_9569_inst flow-through 
    process(B03_9570) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:XOR_u8_u8_9569_inst:flowthrough inputs: " & " A3_9550 = "& Convert_SLV_To_Hex_String(A3_9550) & " Y03x2_9486 = "& Convert_SLV_To_Hex_String(Y03x2_9486) & " outputs:" & " B03_9570= "  & Convert_SLV_To_Hex_String(B03_9570));
      --
    end process; 
    -- binary operator XOR_u8_u8_9569_inst
    process(A3_9550, Y03x2_9486) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(A3_9550, Y03x2_9486, tmp_var);
      B03_9570 <= tmp_var; -- 
    end process;
    -- logger for split-operator XOR_u8_u8_9574_inst flow-through 
    process(B10_9575) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:XOR_u8_u8_9574_inst:flowthrough inputs: " & " A0_9535 = "& Convert_SLV_To_Hex_String(A0_9535) & " Y10x2_9489 = "& Convert_SLV_To_Hex_String(Y10x2_9489) & " outputs:" & " B10_9575= "  & Convert_SLV_To_Hex_String(B10_9575));
      --
    end process; 
    -- binary operator XOR_u8_u8_9574_inst
    process(A0_9535, Y10x2_9489) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(A0_9535, Y10x2_9489, tmp_var);
      B10_9575 <= tmp_var; -- 
    end process;
    -- logger for split-operator XOR_u8_u8_9579_inst flow-through 
    process(B11_9580) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:XOR_u8_u8_9579_inst:flowthrough inputs: " & " A1_9540 = "& Convert_SLV_To_Hex_String(A1_9540) & " Y11x2_9492 = "& Convert_SLV_To_Hex_String(Y11x2_9492) & " outputs:" & " B11_9580= "  & Convert_SLV_To_Hex_String(B11_9580));
      --
    end process; 
    -- binary operator XOR_u8_u8_9579_inst
    process(A1_9540, Y11x2_9492) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(A1_9540, Y11x2_9492, tmp_var);
      B11_9580 <= tmp_var; -- 
    end process;
    -- logger for split-operator XOR_u8_u8_9584_inst flow-through 
    process(B12_9585) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:XOR_u8_u8_9584_inst:flowthrough inputs: " & " A2_9545 = "& Convert_SLV_To_Hex_String(A2_9545) & " Y12x2_9495 = "& Convert_SLV_To_Hex_String(Y12x2_9495) & " outputs:" & " B12_9585= "  & Convert_SLV_To_Hex_String(B12_9585));
      --
    end process; 
    -- binary operator XOR_u8_u8_9584_inst
    process(A2_9545, Y12x2_9495) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(A2_9545, Y12x2_9495, tmp_var);
      B12_9585 <= tmp_var; -- 
    end process;
    -- logger for split-operator XOR_u8_u8_9589_inst flow-through 
    process(B13_9590) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:XOR_u8_u8_9589_inst:flowthrough inputs: " & " A3_9550 = "& Convert_SLV_To_Hex_String(A3_9550) & " Y13x2_9498 = "& Convert_SLV_To_Hex_String(Y13x2_9498) & " outputs:" & " B13_9590= "  & Convert_SLV_To_Hex_String(B13_9590));
      --
    end process; 
    -- binary operator XOR_u8_u8_9589_inst
    process(A3_9550, Y13x2_9498) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(A3_9550, Y13x2_9498, tmp_var);
      B13_9590 <= tmp_var; -- 
    end process;
    -- logger for split-operator XOR_u8_u8_9594_inst flow-through 
    process(XOR_u8_u8_9594_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:XOR_u8_u8_9594_inst:flowthrough inputs: " & " B00_9555 = "& Convert_SLV_To_Hex_String(B00_9555) & " IS00_9290 = "& Convert_SLV_To_Hex_String(IS00_9290) & " outputs:" & " XOR_u8_u8_9594_wire= "  & Convert_SLV_To_Hex_String(XOR_u8_u8_9594_wire));
      --
    end process; 
    -- binary operator XOR_u8_u8_9594_inst
    process(B00_9555, IS00_9290) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(B00_9555, IS00_9290, tmp_var);
      XOR_u8_u8_9594_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator XOR_u8_u8_9597_inst flow-through 
    process(XOR_u8_u8_9597_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:XOR_u8_u8_9597_inst:flowthrough inputs: " & " IS00x2_9353 = "& Convert_SLV_To_Hex_String(IS00x2_9353) & " IS01x2_9356 = "& Convert_SLV_To_Hex_String(IS01x2_9356) & " outputs:" & " XOR_u8_u8_9597_wire= "  & Convert_SLV_To_Hex_String(XOR_u8_u8_9597_wire));
      --
    end process; 
    -- binary operator XOR_u8_u8_9597_inst
    process(IS00x2_9353, IS01x2_9356) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(IS00x2_9353, IS01x2_9356, tmp_var);
      XOR_u8_u8_9597_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator XOR_u8_u8_9598_inst flow-through 
    process(IMX00_9599) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:XOR_u8_u8_9598_inst:flowthrough inputs: " & " XOR_u8_u8_9594_wire = "& Convert_SLV_To_Hex_String(XOR_u8_u8_9594_wire) & " XOR_u8_u8_9597_wire = "& Convert_SLV_To_Hex_String(XOR_u8_u8_9597_wire) & " outputs:" & " IMX00_9599= "  & Convert_SLV_To_Hex_String(IMX00_9599));
      --
    end process; 
    -- binary operator XOR_u8_u8_9598_inst
    process(XOR_u8_u8_9594_wire, XOR_u8_u8_9597_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(XOR_u8_u8_9594_wire, XOR_u8_u8_9597_wire, tmp_var);
      IMX00_9599 <= tmp_var; -- 
    end process;
    -- logger for split-operator XOR_u8_u8_9603_inst flow-through 
    process(XOR_u8_u8_9603_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:XOR_u8_u8_9603_inst:flowthrough inputs: " & " B10_9575 = "& Convert_SLV_To_Hex_String(B10_9575) & " IS01_9294 = "& Convert_SLV_To_Hex_String(IS01_9294) & " outputs:" & " XOR_u8_u8_9603_wire= "  & Convert_SLV_To_Hex_String(XOR_u8_u8_9603_wire));
      --
    end process; 
    -- binary operator XOR_u8_u8_9603_inst
    process(B10_9575, IS01_9294) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(B10_9575, IS01_9294, tmp_var);
      XOR_u8_u8_9603_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator XOR_u8_u8_9606_inst flow-through 
    process(XOR_u8_u8_9606_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:XOR_u8_u8_9606_inst:flowthrough inputs: " & " IS01x2_9356 = "& Convert_SLV_To_Hex_String(IS01x2_9356) & " IS02x2_9359 = "& Convert_SLV_To_Hex_String(IS02x2_9359) & " outputs:" & " XOR_u8_u8_9606_wire= "  & Convert_SLV_To_Hex_String(XOR_u8_u8_9606_wire));
      --
    end process; 
    -- binary operator XOR_u8_u8_9606_inst
    process(IS01x2_9356, IS02x2_9359) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(IS01x2_9356, IS02x2_9359, tmp_var);
      XOR_u8_u8_9606_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator XOR_u8_u8_9607_inst flow-through 
    process(IMX01_9608) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:XOR_u8_u8_9607_inst:flowthrough inputs: " & " XOR_u8_u8_9603_wire = "& Convert_SLV_To_Hex_String(XOR_u8_u8_9603_wire) & " XOR_u8_u8_9606_wire = "& Convert_SLV_To_Hex_String(XOR_u8_u8_9606_wire) & " outputs:" & " IMX01_9608= "  & Convert_SLV_To_Hex_String(IMX01_9608));
      --
    end process; 
    -- binary operator XOR_u8_u8_9607_inst
    process(XOR_u8_u8_9603_wire, XOR_u8_u8_9606_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(XOR_u8_u8_9603_wire, XOR_u8_u8_9606_wire, tmp_var);
      IMX01_9608 <= tmp_var; -- 
    end process;
    -- logger for split-operator XOR_u8_u8_9612_inst flow-through 
    process(XOR_u8_u8_9612_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:XOR_u8_u8_9612_inst:flowthrough inputs: " & " B00_9555 = "& Convert_SLV_To_Hex_String(B00_9555) & " IS02_9298 = "& Convert_SLV_To_Hex_String(IS02_9298) & " outputs:" & " XOR_u8_u8_9612_wire= "  & Convert_SLV_To_Hex_String(XOR_u8_u8_9612_wire));
      --
    end process; 
    -- binary operator XOR_u8_u8_9612_inst
    process(B00_9555, IS02_9298) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(B00_9555, IS02_9298, tmp_var);
      XOR_u8_u8_9612_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator XOR_u8_u8_9615_inst flow-through 
    process(XOR_u8_u8_9615_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:XOR_u8_u8_9615_inst:flowthrough inputs: " & " IS02x2_9359 = "& Convert_SLV_To_Hex_String(IS02x2_9359) & " IS03x2_9362 = "& Convert_SLV_To_Hex_String(IS03x2_9362) & " outputs:" & " XOR_u8_u8_9615_wire= "  & Convert_SLV_To_Hex_String(XOR_u8_u8_9615_wire));
      --
    end process; 
    -- binary operator XOR_u8_u8_9615_inst
    process(IS02x2_9359, IS03x2_9362) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(IS02x2_9359, IS03x2_9362, tmp_var);
      XOR_u8_u8_9615_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator XOR_u8_u8_9616_inst flow-through 
    process(IMX02_9617) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:XOR_u8_u8_9616_inst:flowthrough inputs: " & " XOR_u8_u8_9612_wire = "& Convert_SLV_To_Hex_String(XOR_u8_u8_9612_wire) & " XOR_u8_u8_9615_wire = "& Convert_SLV_To_Hex_String(XOR_u8_u8_9615_wire) & " outputs:" & " IMX02_9617= "  & Convert_SLV_To_Hex_String(IMX02_9617));
      --
    end process; 
    -- binary operator XOR_u8_u8_9616_inst
    process(XOR_u8_u8_9612_wire, XOR_u8_u8_9615_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(XOR_u8_u8_9612_wire, XOR_u8_u8_9615_wire, tmp_var);
      IMX02_9617 <= tmp_var; -- 
    end process;
    -- logger for split-operator XOR_u8_u8_9621_inst flow-through 
    process(XOR_u8_u8_9621_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:XOR_u8_u8_9621_inst:flowthrough inputs: " & " B10_9575 = "& Convert_SLV_To_Hex_String(B10_9575) & " IS03_9302 = "& Convert_SLV_To_Hex_String(IS03_9302) & " outputs:" & " XOR_u8_u8_9621_wire= "  & Convert_SLV_To_Hex_String(XOR_u8_u8_9621_wire));
      --
    end process; 
    -- binary operator XOR_u8_u8_9621_inst
    process(B10_9575, IS03_9302) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(B10_9575, IS03_9302, tmp_var);
      XOR_u8_u8_9621_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator XOR_u8_u8_9624_inst flow-through 
    process(XOR_u8_u8_9624_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:XOR_u8_u8_9624_inst:flowthrough inputs: " & " IS03x2_9362 = "& Convert_SLV_To_Hex_String(IS03x2_9362) & " IS00x2_9353 = "& Convert_SLV_To_Hex_String(IS00x2_9353) & " outputs:" & " XOR_u8_u8_9624_wire= "  & Convert_SLV_To_Hex_String(XOR_u8_u8_9624_wire));
      --
    end process; 
    -- binary operator XOR_u8_u8_9624_inst
    process(IS03x2_9362, IS00x2_9353) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(IS03x2_9362, IS00x2_9353, tmp_var);
      XOR_u8_u8_9624_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator XOR_u8_u8_9625_inst flow-through 
    process(IMX03_9626) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:XOR_u8_u8_9625_inst:flowthrough inputs: " & " XOR_u8_u8_9621_wire = "& Convert_SLV_To_Hex_String(XOR_u8_u8_9621_wire) & " XOR_u8_u8_9624_wire = "& Convert_SLV_To_Hex_String(XOR_u8_u8_9624_wire) & " outputs:" & " IMX03_9626= "  & Convert_SLV_To_Hex_String(IMX03_9626));
      --
    end process; 
    -- binary operator XOR_u8_u8_9625_inst
    process(XOR_u8_u8_9621_wire, XOR_u8_u8_9624_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(XOR_u8_u8_9621_wire, XOR_u8_u8_9624_wire, tmp_var);
      IMX03_9626 <= tmp_var; -- 
    end process;
    -- logger for split-operator XOR_u8_u8_9630_inst flow-through 
    process(XOR_u8_u8_9630_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:XOR_u8_u8_9630_inst:flowthrough inputs: " & " B01_9560 = "& Convert_SLV_To_Hex_String(B01_9560) & " IS04_9306 = "& Convert_SLV_To_Hex_String(IS04_9306) & " outputs:" & " XOR_u8_u8_9630_wire= "  & Convert_SLV_To_Hex_String(XOR_u8_u8_9630_wire));
      --
    end process; 
    -- binary operator XOR_u8_u8_9630_inst
    process(B01_9560, IS04_9306) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(B01_9560, IS04_9306, tmp_var);
      XOR_u8_u8_9630_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator XOR_u8_u8_9633_inst flow-through 
    process(XOR_u8_u8_9633_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:XOR_u8_u8_9633_inst:flowthrough inputs: " & " IS04x2_9365 = "& Convert_SLV_To_Hex_String(IS04x2_9365) & " IS05x2_9368 = "& Convert_SLV_To_Hex_String(IS05x2_9368) & " outputs:" & " XOR_u8_u8_9633_wire= "  & Convert_SLV_To_Hex_String(XOR_u8_u8_9633_wire));
      --
    end process; 
    -- binary operator XOR_u8_u8_9633_inst
    process(IS04x2_9365, IS05x2_9368) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(IS04x2_9365, IS05x2_9368, tmp_var);
      XOR_u8_u8_9633_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator XOR_u8_u8_9634_inst flow-through 
    process(IMX04_9635) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:XOR_u8_u8_9634_inst:flowthrough inputs: " & " XOR_u8_u8_9630_wire = "& Convert_SLV_To_Hex_String(XOR_u8_u8_9630_wire) & " XOR_u8_u8_9633_wire = "& Convert_SLV_To_Hex_String(XOR_u8_u8_9633_wire) & " outputs:" & " IMX04_9635= "  & Convert_SLV_To_Hex_String(IMX04_9635));
      --
    end process; 
    -- binary operator XOR_u8_u8_9634_inst
    process(XOR_u8_u8_9630_wire, XOR_u8_u8_9633_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(XOR_u8_u8_9630_wire, XOR_u8_u8_9633_wire, tmp_var);
      IMX04_9635 <= tmp_var; -- 
    end process;
    -- logger for split-operator XOR_u8_u8_9639_inst flow-through 
    process(XOR_u8_u8_9639_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:XOR_u8_u8_9639_inst:flowthrough inputs: " & " B11_9580 = "& Convert_SLV_To_Hex_String(B11_9580) & " IS05_9310 = "& Convert_SLV_To_Hex_String(IS05_9310) & " outputs:" & " XOR_u8_u8_9639_wire= "  & Convert_SLV_To_Hex_String(XOR_u8_u8_9639_wire));
      --
    end process; 
    -- binary operator XOR_u8_u8_9639_inst
    process(B11_9580, IS05_9310) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(B11_9580, IS05_9310, tmp_var);
      XOR_u8_u8_9639_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator XOR_u8_u8_9642_inst flow-through 
    process(XOR_u8_u8_9642_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:XOR_u8_u8_9642_inst:flowthrough inputs: " & " IS05x2_9368 = "& Convert_SLV_To_Hex_String(IS05x2_9368) & " IS06x2_9371 = "& Convert_SLV_To_Hex_String(IS06x2_9371) & " outputs:" & " XOR_u8_u8_9642_wire= "  & Convert_SLV_To_Hex_String(XOR_u8_u8_9642_wire));
      --
    end process; 
    -- binary operator XOR_u8_u8_9642_inst
    process(IS05x2_9368, IS06x2_9371) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(IS05x2_9368, IS06x2_9371, tmp_var);
      XOR_u8_u8_9642_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator XOR_u8_u8_9643_inst flow-through 
    process(IMX05_9644) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:XOR_u8_u8_9643_inst:flowthrough inputs: " & " XOR_u8_u8_9639_wire = "& Convert_SLV_To_Hex_String(XOR_u8_u8_9639_wire) & " XOR_u8_u8_9642_wire = "& Convert_SLV_To_Hex_String(XOR_u8_u8_9642_wire) & " outputs:" & " IMX05_9644= "  & Convert_SLV_To_Hex_String(IMX05_9644));
      --
    end process; 
    -- binary operator XOR_u8_u8_9643_inst
    process(XOR_u8_u8_9639_wire, XOR_u8_u8_9642_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(XOR_u8_u8_9639_wire, XOR_u8_u8_9642_wire, tmp_var);
      IMX05_9644 <= tmp_var; -- 
    end process;
    -- logger for split-operator XOR_u8_u8_9648_inst flow-through 
    process(XOR_u8_u8_9648_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:XOR_u8_u8_9648_inst:flowthrough inputs: " & " B01_9560 = "& Convert_SLV_To_Hex_String(B01_9560) & " IS06_9314 = "& Convert_SLV_To_Hex_String(IS06_9314) & " outputs:" & " XOR_u8_u8_9648_wire= "  & Convert_SLV_To_Hex_String(XOR_u8_u8_9648_wire));
      --
    end process; 
    -- binary operator XOR_u8_u8_9648_inst
    process(B01_9560, IS06_9314) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(B01_9560, IS06_9314, tmp_var);
      XOR_u8_u8_9648_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator XOR_u8_u8_9651_inst flow-through 
    process(XOR_u8_u8_9651_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:XOR_u8_u8_9651_inst:flowthrough inputs: " & " IS06x2_9371 = "& Convert_SLV_To_Hex_String(IS06x2_9371) & " IS07x2_9374 = "& Convert_SLV_To_Hex_String(IS07x2_9374) & " outputs:" & " XOR_u8_u8_9651_wire= "  & Convert_SLV_To_Hex_String(XOR_u8_u8_9651_wire));
      --
    end process; 
    -- binary operator XOR_u8_u8_9651_inst
    process(IS06x2_9371, IS07x2_9374) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(IS06x2_9371, IS07x2_9374, tmp_var);
      XOR_u8_u8_9651_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator XOR_u8_u8_9652_inst flow-through 
    process(IMX06_9653) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:XOR_u8_u8_9652_inst:flowthrough inputs: " & " XOR_u8_u8_9648_wire = "& Convert_SLV_To_Hex_String(XOR_u8_u8_9648_wire) & " XOR_u8_u8_9651_wire = "& Convert_SLV_To_Hex_String(XOR_u8_u8_9651_wire) & " outputs:" & " IMX06_9653= "  & Convert_SLV_To_Hex_String(IMX06_9653));
      --
    end process; 
    -- binary operator XOR_u8_u8_9652_inst
    process(XOR_u8_u8_9648_wire, XOR_u8_u8_9651_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(XOR_u8_u8_9648_wire, XOR_u8_u8_9651_wire, tmp_var);
      IMX06_9653 <= tmp_var; -- 
    end process;
    -- logger for split-operator XOR_u8_u8_9657_inst flow-through 
    process(XOR_u8_u8_9657_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:XOR_u8_u8_9657_inst:flowthrough inputs: " & " B11_9580 = "& Convert_SLV_To_Hex_String(B11_9580) & " IS07_9318 = "& Convert_SLV_To_Hex_String(IS07_9318) & " outputs:" & " XOR_u8_u8_9657_wire= "  & Convert_SLV_To_Hex_String(XOR_u8_u8_9657_wire));
      --
    end process; 
    -- binary operator XOR_u8_u8_9657_inst
    process(B11_9580, IS07_9318) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(B11_9580, IS07_9318, tmp_var);
      XOR_u8_u8_9657_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator XOR_u8_u8_9660_inst flow-through 
    process(XOR_u8_u8_9660_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:XOR_u8_u8_9660_inst:flowthrough inputs: " & " IS07x2_9374 = "& Convert_SLV_To_Hex_String(IS07x2_9374) & " IS04x2_9365 = "& Convert_SLV_To_Hex_String(IS04x2_9365) & " outputs:" & " XOR_u8_u8_9660_wire= "  & Convert_SLV_To_Hex_String(XOR_u8_u8_9660_wire));
      --
    end process; 
    -- binary operator XOR_u8_u8_9660_inst
    process(IS07x2_9374, IS04x2_9365) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(IS07x2_9374, IS04x2_9365, tmp_var);
      XOR_u8_u8_9660_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator XOR_u8_u8_9661_inst flow-through 
    process(IMX07_9662) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:XOR_u8_u8_9661_inst:flowthrough inputs: " & " XOR_u8_u8_9657_wire = "& Convert_SLV_To_Hex_String(XOR_u8_u8_9657_wire) & " XOR_u8_u8_9660_wire = "& Convert_SLV_To_Hex_String(XOR_u8_u8_9660_wire) & " outputs:" & " IMX07_9662= "  & Convert_SLV_To_Hex_String(IMX07_9662));
      --
    end process; 
    -- binary operator XOR_u8_u8_9661_inst
    process(XOR_u8_u8_9657_wire, XOR_u8_u8_9660_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(XOR_u8_u8_9657_wire, XOR_u8_u8_9660_wire, tmp_var);
      IMX07_9662 <= tmp_var; -- 
    end process;
    -- logger for split-operator XOR_u8_u8_9666_inst flow-through 
    process(XOR_u8_u8_9666_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:XOR_u8_u8_9666_inst:flowthrough inputs: " & " B02_9565 = "& Convert_SLV_To_Hex_String(B02_9565) & " IS08_9322 = "& Convert_SLV_To_Hex_String(IS08_9322) & " outputs:" & " XOR_u8_u8_9666_wire= "  & Convert_SLV_To_Hex_String(XOR_u8_u8_9666_wire));
      --
    end process; 
    -- binary operator XOR_u8_u8_9666_inst
    process(B02_9565, IS08_9322) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(B02_9565, IS08_9322, tmp_var);
      XOR_u8_u8_9666_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator XOR_u8_u8_9669_inst flow-through 
    process(XOR_u8_u8_9669_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:XOR_u8_u8_9669_inst:flowthrough inputs: " & " IS08x2_9377 = "& Convert_SLV_To_Hex_String(IS08x2_9377) & " IS09x2_9380 = "& Convert_SLV_To_Hex_String(IS09x2_9380) & " outputs:" & " XOR_u8_u8_9669_wire= "  & Convert_SLV_To_Hex_String(XOR_u8_u8_9669_wire));
      --
    end process; 
    -- binary operator XOR_u8_u8_9669_inst
    process(IS08x2_9377, IS09x2_9380) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(IS08x2_9377, IS09x2_9380, tmp_var);
      XOR_u8_u8_9669_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator XOR_u8_u8_9670_inst flow-through 
    process(IMX08_9671) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:XOR_u8_u8_9670_inst:flowthrough inputs: " & " XOR_u8_u8_9666_wire = "& Convert_SLV_To_Hex_String(XOR_u8_u8_9666_wire) & " XOR_u8_u8_9669_wire = "& Convert_SLV_To_Hex_String(XOR_u8_u8_9669_wire) & " outputs:" & " IMX08_9671= "  & Convert_SLV_To_Hex_String(IMX08_9671));
      --
    end process; 
    -- binary operator XOR_u8_u8_9670_inst
    process(XOR_u8_u8_9666_wire, XOR_u8_u8_9669_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(XOR_u8_u8_9666_wire, XOR_u8_u8_9669_wire, tmp_var);
      IMX08_9671 <= tmp_var; -- 
    end process;
    -- logger for split-operator XOR_u8_u8_9675_inst flow-through 
    process(XOR_u8_u8_9675_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:XOR_u8_u8_9675_inst:flowthrough inputs: " & " B12_9585 = "& Convert_SLV_To_Hex_String(B12_9585) & " IS09_9326 = "& Convert_SLV_To_Hex_String(IS09_9326) & " outputs:" & " XOR_u8_u8_9675_wire= "  & Convert_SLV_To_Hex_String(XOR_u8_u8_9675_wire));
      --
    end process; 
    -- binary operator XOR_u8_u8_9675_inst
    process(B12_9585, IS09_9326) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(B12_9585, IS09_9326, tmp_var);
      XOR_u8_u8_9675_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator XOR_u8_u8_9678_inst flow-through 
    process(XOR_u8_u8_9678_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:XOR_u8_u8_9678_inst:flowthrough inputs: " & " IS09x2_9380 = "& Convert_SLV_To_Hex_String(IS09x2_9380) & " IS10x2_9383 = "& Convert_SLV_To_Hex_String(IS10x2_9383) & " outputs:" & " XOR_u8_u8_9678_wire= "  & Convert_SLV_To_Hex_String(XOR_u8_u8_9678_wire));
      --
    end process; 
    -- binary operator XOR_u8_u8_9678_inst
    process(IS09x2_9380, IS10x2_9383) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(IS09x2_9380, IS10x2_9383, tmp_var);
      XOR_u8_u8_9678_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator XOR_u8_u8_9679_inst flow-through 
    process(IMX09_9680) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:XOR_u8_u8_9679_inst:flowthrough inputs: " & " XOR_u8_u8_9675_wire = "& Convert_SLV_To_Hex_String(XOR_u8_u8_9675_wire) & " XOR_u8_u8_9678_wire = "& Convert_SLV_To_Hex_String(XOR_u8_u8_9678_wire) & " outputs:" & " IMX09_9680= "  & Convert_SLV_To_Hex_String(IMX09_9680));
      --
    end process; 
    -- binary operator XOR_u8_u8_9679_inst
    process(XOR_u8_u8_9675_wire, XOR_u8_u8_9678_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(XOR_u8_u8_9675_wire, XOR_u8_u8_9678_wire, tmp_var);
      IMX09_9680 <= tmp_var; -- 
    end process;
    -- logger for split-operator XOR_u8_u8_9684_inst flow-through 
    process(XOR_u8_u8_9684_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:XOR_u8_u8_9684_inst:flowthrough inputs: " & " B02_9565 = "& Convert_SLV_To_Hex_String(B02_9565) & " IS10_9330 = "& Convert_SLV_To_Hex_String(IS10_9330) & " outputs:" & " XOR_u8_u8_9684_wire= "  & Convert_SLV_To_Hex_String(XOR_u8_u8_9684_wire));
      --
    end process; 
    -- binary operator XOR_u8_u8_9684_inst
    process(B02_9565, IS10_9330) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(B02_9565, IS10_9330, tmp_var);
      XOR_u8_u8_9684_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator XOR_u8_u8_9687_inst flow-through 
    process(XOR_u8_u8_9687_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:XOR_u8_u8_9687_inst:flowthrough inputs: " & " IS10x2_9383 = "& Convert_SLV_To_Hex_String(IS10x2_9383) & " IS11x2_9386 = "& Convert_SLV_To_Hex_String(IS11x2_9386) & " outputs:" & " XOR_u8_u8_9687_wire= "  & Convert_SLV_To_Hex_String(XOR_u8_u8_9687_wire));
      --
    end process; 
    -- binary operator XOR_u8_u8_9687_inst
    process(IS10x2_9383, IS11x2_9386) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(IS10x2_9383, IS11x2_9386, tmp_var);
      XOR_u8_u8_9687_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator XOR_u8_u8_9688_inst flow-through 
    process(IMX10_9689) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:XOR_u8_u8_9688_inst:flowthrough inputs: " & " XOR_u8_u8_9684_wire = "& Convert_SLV_To_Hex_String(XOR_u8_u8_9684_wire) & " XOR_u8_u8_9687_wire = "& Convert_SLV_To_Hex_String(XOR_u8_u8_9687_wire) & " outputs:" & " IMX10_9689= "  & Convert_SLV_To_Hex_String(IMX10_9689));
      --
    end process; 
    -- binary operator XOR_u8_u8_9688_inst
    process(XOR_u8_u8_9684_wire, XOR_u8_u8_9687_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(XOR_u8_u8_9684_wire, XOR_u8_u8_9687_wire, tmp_var);
      IMX10_9689 <= tmp_var; -- 
    end process;
    -- logger for split-operator XOR_u8_u8_9693_inst flow-through 
    process(XOR_u8_u8_9693_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:XOR_u8_u8_9693_inst:flowthrough inputs: " & " B12_9585 = "& Convert_SLV_To_Hex_String(B12_9585) & " IS11_9334 = "& Convert_SLV_To_Hex_String(IS11_9334) & " outputs:" & " XOR_u8_u8_9693_wire= "  & Convert_SLV_To_Hex_String(XOR_u8_u8_9693_wire));
      --
    end process; 
    -- binary operator XOR_u8_u8_9693_inst
    process(B12_9585, IS11_9334) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(B12_9585, IS11_9334, tmp_var);
      XOR_u8_u8_9693_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator XOR_u8_u8_9696_inst flow-through 
    process(XOR_u8_u8_9696_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:XOR_u8_u8_9696_inst:flowthrough inputs: " & " IS11x2_9386 = "& Convert_SLV_To_Hex_String(IS11x2_9386) & " IS08x2_9377 = "& Convert_SLV_To_Hex_String(IS08x2_9377) & " outputs:" & " XOR_u8_u8_9696_wire= "  & Convert_SLV_To_Hex_String(XOR_u8_u8_9696_wire));
      --
    end process; 
    -- binary operator XOR_u8_u8_9696_inst
    process(IS11x2_9386, IS08x2_9377) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(IS11x2_9386, IS08x2_9377, tmp_var);
      XOR_u8_u8_9696_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator XOR_u8_u8_9697_inst flow-through 
    process(IMX11_9698) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:XOR_u8_u8_9697_inst:flowthrough inputs: " & " XOR_u8_u8_9693_wire = "& Convert_SLV_To_Hex_String(XOR_u8_u8_9693_wire) & " XOR_u8_u8_9696_wire = "& Convert_SLV_To_Hex_String(XOR_u8_u8_9696_wire) & " outputs:" & " IMX11_9698= "  & Convert_SLV_To_Hex_String(IMX11_9698));
      --
    end process; 
    -- binary operator XOR_u8_u8_9697_inst
    process(XOR_u8_u8_9693_wire, XOR_u8_u8_9696_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(XOR_u8_u8_9693_wire, XOR_u8_u8_9696_wire, tmp_var);
      IMX11_9698 <= tmp_var; -- 
    end process;
    -- logger for split-operator XOR_u8_u8_9702_inst flow-through 
    process(XOR_u8_u8_9702_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:XOR_u8_u8_9702_inst:flowthrough inputs: " & " B03_9570 = "& Convert_SLV_To_Hex_String(B03_9570) & " IS12_9338 = "& Convert_SLV_To_Hex_String(IS12_9338) & " outputs:" & " XOR_u8_u8_9702_wire= "  & Convert_SLV_To_Hex_String(XOR_u8_u8_9702_wire));
      --
    end process; 
    -- binary operator XOR_u8_u8_9702_inst
    process(B03_9570, IS12_9338) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(B03_9570, IS12_9338, tmp_var);
      XOR_u8_u8_9702_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator XOR_u8_u8_9705_inst flow-through 
    process(XOR_u8_u8_9705_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:XOR_u8_u8_9705_inst:flowthrough inputs: " & " IS12x2_9389 = "& Convert_SLV_To_Hex_String(IS12x2_9389) & " IS13x2_9392 = "& Convert_SLV_To_Hex_String(IS13x2_9392) & " outputs:" & " XOR_u8_u8_9705_wire= "  & Convert_SLV_To_Hex_String(XOR_u8_u8_9705_wire));
      --
    end process; 
    -- binary operator XOR_u8_u8_9705_inst
    process(IS12x2_9389, IS13x2_9392) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(IS12x2_9389, IS13x2_9392, tmp_var);
      XOR_u8_u8_9705_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator XOR_u8_u8_9706_inst flow-through 
    process(IMX12_9707) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:XOR_u8_u8_9706_inst:flowthrough inputs: " & " XOR_u8_u8_9702_wire = "& Convert_SLV_To_Hex_String(XOR_u8_u8_9702_wire) & " XOR_u8_u8_9705_wire = "& Convert_SLV_To_Hex_String(XOR_u8_u8_9705_wire) & " outputs:" & " IMX12_9707= "  & Convert_SLV_To_Hex_String(IMX12_9707));
      --
    end process; 
    -- binary operator XOR_u8_u8_9706_inst
    process(XOR_u8_u8_9702_wire, XOR_u8_u8_9705_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(XOR_u8_u8_9702_wire, XOR_u8_u8_9705_wire, tmp_var);
      IMX12_9707 <= tmp_var; -- 
    end process;
    -- logger for split-operator XOR_u8_u8_9711_inst flow-through 
    process(XOR_u8_u8_9711_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:XOR_u8_u8_9711_inst:flowthrough inputs: " & " B13_9590 = "& Convert_SLV_To_Hex_String(B13_9590) & " IS13_9342 = "& Convert_SLV_To_Hex_String(IS13_9342) & " outputs:" & " XOR_u8_u8_9711_wire= "  & Convert_SLV_To_Hex_String(XOR_u8_u8_9711_wire));
      --
    end process; 
    -- binary operator XOR_u8_u8_9711_inst
    process(B13_9590, IS13_9342) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(B13_9590, IS13_9342, tmp_var);
      XOR_u8_u8_9711_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator XOR_u8_u8_9714_inst flow-through 
    process(XOR_u8_u8_9714_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:XOR_u8_u8_9714_inst:flowthrough inputs: " & " IS13x2_9392 = "& Convert_SLV_To_Hex_String(IS13x2_9392) & " IS14x2_9395 = "& Convert_SLV_To_Hex_String(IS14x2_9395) & " outputs:" & " XOR_u8_u8_9714_wire= "  & Convert_SLV_To_Hex_String(XOR_u8_u8_9714_wire));
      --
    end process; 
    -- binary operator XOR_u8_u8_9714_inst
    process(IS13x2_9392, IS14x2_9395) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(IS13x2_9392, IS14x2_9395, tmp_var);
      XOR_u8_u8_9714_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator XOR_u8_u8_9715_inst flow-through 
    process(IMX13_9716) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:XOR_u8_u8_9715_inst:flowthrough inputs: " & " XOR_u8_u8_9711_wire = "& Convert_SLV_To_Hex_String(XOR_u8_u8_9711_wire) & " XOR_u8_u8_9714_wire = "& Convert_SLV_To_Hex_String(XOR_u8_u8_9714_wire) & " outputs:" & " IMX13_9716= "  & Convert_SLV_To_Hex_String(IMX13_9716));
      --
    end process; 
    -- binary operator XOR_u8_u8_9715_inst
    process(XOR_u8_u8_9711_wire, XOR_u8_u8_9714_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(XOR_u8_u8_9711_wire, XOR_u8_u8_9714_wire, tmp_var);
      IMX13_9716 <= tmp_var; -- 
    end process;
    -- logger for split-operator XOR_u8_u8_9720_inst flow-through 
    process(XOR_u8_u8_9720_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:XOR_u8_u8_9720_inst:flowthrough inputs: " & " B03_9570 = "& Convert_SLV_To_Hex_String(B03_9570) & " IS14_9346 = "& Convert_SLV_To_Hex_String(IS14_9346) & " outputs:" & " XOR_u8_u8_9720_wire= "  & Convert_SLV_To_Hex_String(XOR_u8_u8_9720_wire));
      --
    end process; 
    -- binary operator XOR_u8_u8_9720_inst
    process(B03_9570, IS14_9346) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(B03_9570, IS14_9346, tmp_var);
      XOR_u8_u8_9720_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator XOR_u8_u8_9723_inst flow-through 
    process(XOR_u8_u8_9723_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:XOR_u8_u8_9723_inst:flowthrough inputs: " & " IS14x2_9395 = "& Convert_SLV_To_Hex_String(IS14x2_9395) & " IS15x2_9398 = "& Convert_SLV_To_Hex_String(IS15x2_9398) & " outputs:" & " XOR_u8_u8_9723_wire= "  & Convert_SLV_To_Hex_String(XOR_u8_u8_9723_wire));
      --
    end process; 
    -- binary operator XOR_u8_u8_9723_inst
    process(IS14x2_9395, IS15x2_9398) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(IS14x2_9395, IS15x2_9398, tmp_var);
      XOR_u8_u8_9723_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator XOR_u8_u8_9724_inst flow-through 
    process(IMX14_9725) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:XOR_u8_u8_9724_inst:flowthrough inputs: " & " XOR_u8_u8_9720_wire = "& Convert_SLV_To_Hex_String(XOR_u8_u8_9720_wire) & " XOR_u8_u8_9723_wire = "& Convert_SLV_To_Hex_String(XOR_u8_u8_9723_wire) & " outputs:" & " IMX14_9725= "  & Convert_SLV_To_Hex_String(IMX14_9725));
      --
    end process; 
    -- binary operator XOR_u8_u8_9724_inst
    process(XOR_u8_u8_9720_wire, XOR_u8_u8_9723_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(XOR_u8_u8_9720_wire, XOR_u8_u8_9723_wire, tmp_var);
      IMX14_9725 <= tmp_var; -- 
    end process;
    -- logger for split-operator XOR_u8_u8_9729_inst flow-through 
    process(XOR_u8_u8_9729_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:XOR_u8_u8_9729_inst:flowthrough inputs: " & " B13_9590 = "& Convert_SLV_To_Hex_String(B13_9590) & " IS15_9350 = "& Convert_SLV_To_Hex_String(IS15_9350) & " outputs:" & " XOR_u8_u8_9729_wire= "  & Convert_SLV_To_Hex_String(XOR_u8_u8_9729_wire));
      --
    end process; 
    -- binary operator XOR_u8_u8_9729_inst
    process(B13_9590, IS15_9350) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(B13_9590, IS15_9350, tmp_var);
      XOR_u8_u8_9729_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator XOR_u8_u8_9732_inst flow-through 
    process(XOR_u8_u8_9732_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:XOR_u8_u8_9732_inst:flowthrough inputs: " & " IS15x2_9398 = "& Convert_SLV_To_Hex_String(IS15x2_9398) & " IS12x2_9389 = "& Convert_SLV_To_Hex_String(IS12x2_9389) & " outputs:" & " XOR_u8_u8_9732_wire= "  & Convert_SLV_To_Hex_String(XOR_u8_u8_9732_wire));
      --
    end process; 
    -- binary operator XOR_u8_u8_9732_inst
    process(IS15x2_9398, IS12x2_9389) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(IS15x2_9398, IS12x2_9389, tmp_var);
      XOR_u8_u8_9732_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator XOR_u8_u8_9733_inst flow-through 
    process(IMX15_9734) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:XOR_u8_u8_9733_inst:flowthrough inputs: " & " XOR_u8_u8_9729_wire = "& Convert_SLV_To_Hex_String(XOR_u8_u8_9729_wire) & " XOR_u8_u8_9732_wire = "& Convert_SLV_To_Hex_String(XOR_u8_u8_9732_wire) & " outputs:" & " IMX15_9734= "  & Convert_SLV_To_Hex_String(IMX15_9734));
      --
    end process; 
    -- binary operator XOR_u8_u8_9733_inst
    process(XOR_u8_u8_9729_wire, XOR_u8_u8_9732_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(XOR_u8_u8_9729_wire, XOR_u8_u8_9732_wire, tmp_var);
      IMX15_9734 <= tmp_var; -- 
    end process;
    -- logger for split-operator call_stmt_9353_call flow-through 
    process(IS00x2_9353) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:call_stmt_9353_call:flowthrough inputs: " & " IS00_9290 = "& Convert_SLV_To_Hex_String(IS00_9290) & " outputs:" & " IS00x2_9353= "  & Convert_SLV_To_Hex_String(IS00x2_9353));
      --
    end process; 
    call_inst_11762: MUL2_Volatile port map(mul_in => IS00_9290, mul_out => IS00x2_9353, clk => clk, reset => reset); 
    -- logger for split-operator call_stmt_9356_call flow-through 
    process(IS01x2_9356) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:call_stmt_9356_call:flowthrough inputs: " & " IS01_9294 = "& Convert_SLV_To_Hex_String(IS01_9294) & " outputs:" & " IS01x2_9356= "  & Convert_SLV_To_Hex_String(IS01x2_9356));
      --
    end process; 
    call_inst_11763: MUL2_Volatile port map(mul_in => IS01_9294, mul_out => IS01x2_9356, clk => clk, reset => reset); 
    -- logger for split-operator call_stmt_9359_call flow-through 
    process(IS02x2_9359) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:call_stmt_9359_call:flowthrough inputs: " & " IS02_9298 = "& Convert_SLV_To_Hex_String(IS02_9298) & " outputs:" & " IS02x2_9359= "  & Convert_SLV_To_Hex_String(IS02x2_9359));
      --
    end process; 
    call_inst_11764: MUL2_Volatile port map(mul_in => IS02_9298, mul_out => IS02x2_9359, clk => clk, reset => reset); 
    -- logger for split-operator call_stmt_9362_call flow-through 
    process(IS03x2_9362) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:call_stmt_9362_call:flowthrough inputs: " & " IS03_9302 = "& Convert_SLV_To_Hex_String(IS03_9302) & " outputs:" & " IS03x2_9362= "  & Convert_SLV_To_Hex_String(IS03x2_9362));
      --
    end process; 
    call_inst_11765: MUL2_Volatile port map(mul_in => IS03_9302, mul_out => IS03x2_9362, clk => clk, reset => reset); 
    -- logger for split-operator call_stmt_9365_call flow-through 
    process(IS04x2_9365) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:call_stmt_9365_call:flowthrough inputs: " & " IS04_9306 = "& Convert_SLV_To_Hex_String(IS04_9306) & " outputs:" & " IS04x2_9365= "  & Convert_SLV_To_Hex_String(IS04x2_9365));
      --
    end process; 
    call_inst_11766: MUL2_Volatile port map(mul_in => IS04_9306, mul_out => IS04x2_9365, clk => clk, reset => reset); 
    -- logger for split-operator call_stmt_9368_call flow-through 
    process(IS05x2_9368) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:call_stmt_9368_call:flowthrough inputs: " & " IS05_9310 = "& Convert_SLV_To_Hex_String(IS05_9310) & " outputs:" & " IS05x2_9368= "  & Convert_SLV_To_Hex_String(IS05x2_9368));
      --
    end process; 
    call_inst_11767: MUL2_Volatile port map(mul_in => IS05_9310, mul_out => IS05x2_9368, clk => clk, reset => reset); 
    -- logger for split-operator call_stmt_9371_call flow-through 
    process(IS06x2_9371) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:call_stmt_9371_call:flowthrough inputs: " & " IS06_9314 = "& Convert_SLV_To_Hex_String(IS06_9314) & " outputs:" & " IS06x2_9371= "  & Convert_SLV_To_Hex_String(IS06x2_9371));
      --
    end process; 
    call_inst_11768: MUL2_Volatile port map(mul_in => IS06_9314, mul_out => IS06x2_9371, clk => clk, reset => reset); 
    -- logger for split-operator call_stmt_9374_call flow-through 
    process(IS07x2_9374) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:call_stmt_9374_call:flowthrough inputs: " & " IS07_9318 = "& Convert_SLV_To_Hex_String(IS07_9318) & " outputs:" & " IS07x2_9374= "  & Convert_SLV_To_Hex_String(IS07x2_9374));
      --
    end process; 
    call_inst_11769: MUL2_Volatile port map(mul_in => IS07_9318, mul_out => IS07x2_9374, clk => clk, reset => reset); 
    -- logger for split-operator call_stmt_9377_call flow-through 
    process(IS08x2_9377) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:call_stmt_9377_call:flowthrough inputs: " & " IS08_9322 = "& Convert_SLV_To_Hex_String(IS08_9322) & " outputs:" & " IS08x2_9377= "  & Convert_SLV_To_Hex_String(IS08x2_9377));
      --
    end process; 
    call_inst_11770: MUL2_Volatile port map(mul_in => IS08_9322, mul_out => IS08x2_9377, clk => clk, reset => reset); 
    -- logger for split-operator call_stmt_9380_call flow-through 
    process(IS09x2_9380) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:call_stmt_9380_call:flowthrough inputs: " & " IS09_9326 = "& Convert_SLV_To_Hex_String(IS09_9326) & " outputs:" & " IS09x2_9380= "  & Convert_SLV_To_Hex_String(IS09x2_9380));
      --
    end process; 
    call_inst_11771: MUL2_Volatile port map(mul_in => IS09_9326, mul_out => IS09x2_9380, clk => clk, reset => reset); 
    -- logger for split-operator call_stmt_9383_call flow-through 
    process(IS10x2_9383) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:call_stmt_9383_call:flowthrough inputs: " & " IS10_9330 = "& Convert_SLV_To_Hex_String(IS10_9330) & " outputs:" & " IS10x2_9383= "  & Convert_SLV_To_Hex_String(IS10x2_9383));
      --
    end process; 
    call_inst_11772: MUL2_Volatile port map(mul_in => IS10_9330, mul_out => IS10x2_9383, clk => clk, reset => reset); 
    -- logger for split-operator call_stmt_9386_call flow-through 
    process(IS11x2_9386) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:call_stmt_9386_call:flowthrough inputs: " & " IS11_9334 = "& Convert_SLV_To_Hex_String(IS11_9334) & " outputs:" & " IS11x2_9386= "  & Convert_SLV_To_Hex_String(IS11x2_9386));
      --
    end process; 
    call_inst_11773: MUL2_Volatile port map(mul_in => IS11_9334, mul_out => IS11x2_9386, clk => clk, reset => reset); 
    -- logger for split-operator call_stmt_9389_call flow-through 
    process(IS12x2_9389) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:call_stmt_9389_call:flowthrough inputs: " & " IS12_9338 = "& Convert_SLV_To_Hex_String(IS12_9338) & " outputs:" & " IS12x2_9389= "  & Convert_SLV_To_Hex_String(IS12x2_9389));
      --
    end process; 
    call_inst_11774: MUL2_Volatile port map(mul_in => IS12_9338, mul_out => IS12x2_9389, clk => clk, reset => reset); 
    -- logger for split-operator call_stmt_9392_call flow-through 
    process(IS13x2_9392) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:call_stmt_9392_call:flowthrough inputs: " & " IS13_9342 = "& Convert_SLV_To_Hex_String(IS13_9342) & " outputs:" & " IS13x2_9392= "  & Convert_SLV_To_Hex_String(IS13x2_9392));
      --
    end process; 
    call_inst_11775: MUL2_Volatile port map(mul_in => IS13_9342, mul_out => IS13x2_9392, clk => clk, reset => reset); 
    -- logger for split-operator call_stmt_9395_call flow-through 
    process(IS14x2_9395) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:call_stmt_9395_call:flowthrough inputs: " & " IS14_9346 = "& Convert_SLV_To_Hex_String(IS14_9346) & " outputs:" & " IS14x2_9395= "  & Convert_SLV_To_Hex_String(IS14x2_9395));
      --
    end process; 
    call_inst_11776: MUL2_Volatile port map(mul_in => IS14_9346, mul_out => IS14x2_9395, clk => clk, reset => reset); 
    -- logger for split-operator call_stmt_9398_call flow-through 
    process(IS15x2_9398) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:call_stmt_9398_call:flowthrough inputs: " & " IS15_9350 = "& Convert_SLV_To_Hex_String(IS15_9350) & " outputs:" & " IS15x2_9398= "  & Convert_SLV_To_Hex_String(IS15x2_9398));
      --
    end process; 
    call_inst_11777: MUL2_Volatile port map(mul_in => IS15_9350, mul_out => IS15x2_9398, clk => clk, reset => reset); 
    -- logger for split-operator call_stmt_9477_call flow-through 
    process(Y00x2_9477) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:call_stmt_9477_call:flowthrough inputs: " & " Y00_9439 = "& Convert_SLV_To_Hex_String(Y00_9439) & " outputs:" & " Y00x2_9477= "  & Convert_SLV_To_Hex_String(Y00x2_9477));
      --
    end process; 
    call_inst_11798: MUL2_Volatile port map(mul_in => Y00_9439, mul_out => Y00x2_9477, clk => clk, reset => reset); 
    -- logger for split-operator call_stmt_9480_call flow-through 
    process(Y01x2_9480) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:call_stmt_9480_call:flowthrough inputs: " & " Y01_9444 = "& Convert_SLV_To_Hex_String(Y01_9444) & " outputs:" & " Y01x2_9480= "  & Convert_SLV_To_Hex_String(Y01x2_9480));
      --
    end process; 
    call_inst_11799: MUL2_Volatile port map(mul_in => Y01_9444, mul_out => Y01x2_9480, clk => clk, reset => reset); 
    -- logger for split-operator call_stmt_9483_call flow-through 
    process(Y02x2_9483) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:call_stmt_9483_call:flowthrough inputs: " & " Y02_9449 = "& Convert_SLV_To_Hex_String(Y02_9449) & " outputs:" & " Y02x2_9483= "  & Convert_SLV_To_Hex_String(Y02x2_9483));
      --
    end process; 
    call_inst_11800: MUL2_Volatile port map(mul_in => Y02_9449, mul_out => Y02x2_9483, clk => clk, reset => reset); 
    -- logger for split-operator call_stmt_9486_call flow-through 
    process(Y03x2_9486) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:call_stmt_9486_call:flowthrough inputs: " & " Y03_9454 = "& Convert_SLV_To_Hex_String(Y03_9454) & " outputs:" & " Y03x2_9486= "  & Convert_SLV_To_Hex_String(Y03x2_9486));
      --
    end process; 
    call_inst_11801: MUL2_Volatile port map(mul_in => Y03_9454, mul_out => Y03x2_9486, clk => clk, reset => reset); 
    -- logger for split-operator call_stmt_9489_call flow-through 
    process(Y10x2_9489) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:call_stmt_9489_call:flowthrough inputs: " & " Y10_9459 = "& Convert_SLV_To_Hex_String(Y10_9459) & " outputs:" & " Y10x2_9489= "  & Convert_SLV_To_Hex_String(Y10x2_9489));
      --
    end process; 
    call_inst_11802: MUL2_Volatile port map(mul_in => Y10_9459, mul_out => Y10x2_9489, clk => clk, reset => reset); 
    -- logger for split-operator call_stmt_9492_call flow-through 
    process(Y11x2_9492) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:call_stmt_9492_call:flowthrough inputs: " & " Y11_9464 = "& Convert_SLV_To_Hex_String(Y11_9464) & " outputs:" & " Y11x2_9492= "  & Convert_SLV_To_Hex_String(Y11x2_9492));
      --
    end process; 
    call_inst_11803: MUL2_Volatile port map(mul_in => Y11_9464, mul_out => Y11x2_9492, clk => clk, reset => reset); 
    -- logger for split-operator call_stmt_9495_call flow-through 
    process(Y12x2_9495) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:call_stmt_9495_call:flowthrough inputs: " & " Y12_9469 = "& Convert_SLV_To_Hex_String(Y12_9469) & " outputs:" & " Y12x2_9495= "  & Convert_SLV_To_Hex_String(Y12x2_9495));
      --
    end process; 
    call_inst_11804: MUL2_Volatile port map(mul_in => Y12_9469, mul_out => Y12x2_9495, clk => clk, reset => reset); 
    -- logger for split-operator call_stmt_9498_call flow-through 
    process(Y13x2_9498) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:call_stmt_9498_call:flowthrough inputs: " & " Y13_9474 = "& Convert_SLV_To_Hex_String(Y13_9474) & " outputs:" & " Y13x2_9498= "  & Convert_SLV_To_Hex_String(Y13x2_9498));
      --
    end process; 
    call_inst_11805: MUL2_Volatile port map(mul_in => Y13_9474, mul_out => Y13x2_9498, clk => clk, reset => reset); 
    -- logger for split-operator call_stmt_9521_call flow-through 
    process(Z0x2_9521) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:call_stmt_9521_call:flowthrough inputs: " & " Z0_9503 = "& Convert_SLV_To_Hex_String(Z0_9503) & " outputs:" & " Z0x2_9521= "  & Convert_SLV_To_Hex_String(Z0x2_9521));
      --
    end process; 
    call_inst_11810: MUL2_Volatile port map(mul_in => Z0_9503, mul_out => Z0x2_9521, clk => clk, reset => reset); 
    -- logger for split-operator call_stmt_9524_call flow-through 
    process(Z1x2_9524) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:call_stmt_9524_call:flowthrough inputs: " & " Z1_9508 = "& Convert_SLV_To_Hex_String(Z1_9508) & " outputs:" & " Z1x2_9524= "  & Convert_SLV_To_Hex_String(Z1x2_9524));
      --
    end process; 
    call_inst_11811: MUL2_Volatile port map(mul_in => Z1_9508, mul_out => Z1x2_9524, clk => clk, reset => reset); 
    -- logger for split-operator call_stmt_9527_call flow-through 
    process(Z2x2_9527) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:call_stmt_9527_call:flowthrough inputs: " & " Z2_9513 = "& Convert_SLV_To_Hex_String(Z2_9513) & " outputs:" & " Z2x2_9527= "  & Convert_SLV_To_Hex_String(Z2x2_9527));
      --
    end process; 
    call_inst_11812: MUL2_Volatile port map(mul_in => Z2_9513, mul_out => Z2x2_9527, clk => clk, reset => reset); 
    -- logger for split-operator call_stmt_9530_call flow-through 
    process(Z3x2_9530) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:call_stmt_9530_call:flowthrough inputs: " & " Z3_9518 = "& Convert_SLV_To_Hex_String(Z3_9518) & " outputs:" & " Z3x2_9530= "  & Convert_SLV_To_Hex_String(Z3x2_9530));
      --
    end process; 
    call_inst_11813: MUL2_Volatile port map(mul_in => Z3_9518, mul_out => Z3x2_9530, clk => clk, reset => reset); 
    -- logger for split-operator call_stmt_9833_call flow-through 
    process(Sout00_9833) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:call_stmt_9833_call:flowthrough inputs: " & " ISbox_in00_9740 = "& Convert_SLV_To_Hex_String(ISbox_in00_9740) & " outputs:" & " Sout00_9833= "  & Convert_SLV_To_Hex_String(Sout00_9833));
      --
    end process; 
    call_inst_11890: Inv_Sbox_1_Volatile port map(s_in => ISbox_in00_9740, s_out => Sout00_9833, clk => clk, reset => reset); 
    -- logger for split-operator call_stmt_9836_call flow-through 
    process(Sout05_9836) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:call_stmt_9836_call:flowthrough inputs: " & " ISbox_in01_9746 = "& Convert_SLV_To_Hex_String(ISbox_in01_9746) & " outputs:" & " Sout05_9836= "  & Convert_SLV_To_Hex_String(Sout05_9836));
      --
    end process; 
    call_inst_11891: Inv_Sbox_2_Volatile port map(s_in => ISbox_in01_9746, s_out => Sout05_9836, clk => clk, reset => reset); 
    -- logger for split-operator call_stmt_9839_call flow-through 
    process(Sout10_9839) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:call_stmt_9839_call:flowthrough inputs: " & " ISbox_in02_9752 = "& Convert_SLV_To_Hex_String(ISbox_in02_9752) & " outputs:" & " Sout10_9839= "  & Convert_SLV_To_Hex_String(Sout10_9839));
      --
    end process; 
    call_inst_11892: Inv_Sbox_3_Volatile port map(s_in => ISbox_in02_9752, s_out => Sout10_9839, clk => clk, reset => reset); 
    -- logger for split-operator call_stmt_9842_call flow-through 
    process(Sout15_9842) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:call_stmt_9842_call:flowthrough inputs: " & " ISbox_in03_9758 = "& Convert_SLV_To_Hex_String(ISbox_in03_9758) & " outputs:" & " Sout15_9842= "  & Convert_SLV_To_Hex_String(Sout15_9842));
      --
    end process; 
    call_inst_11893: Inv_Sbox_4_Volatile port map(s_in => ISbox_in03_9758, s_out => Sout15_9842, clk => clk, reset => reset); 
    -- logger for split-operator call_stmt_9845_call flow-through 
    process(Sout04_9845) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:call_stmt_9845_call:flowthrough inputs: " & " ISbox_in04_9764 = "& Convert_SLV_To_Hex_String(ISbox_in04_9764) & " outputs:" & " Sout04_9845= "  & Convert_SLV_To_Hex_String(Sout04_9845));
      --
    end process; 
    call_inst_11894: Inv_Sbox_1_Volatile port map(s_in => ISbox_in04_9764, s_out => Sout04_9845, clk => clk, reset => reset); 
    -- logger for split-operator call_stmt_9848_call flow-through 
    process(Sout09_9848) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:call_stmt_9848_call:flowthrough inputs: " & " ISbox_in05_9770 = "& Convert_SLV_To_Hex_String(ISbox_in05_9770) & " outputs:" & " Sout09_9848= "  & Convert_SLV_To_Hex_String(Sout09_9848));
      --
    end process; 
    call_inst_11895: Inv_Sbox_2_Volatile port map(s_in => ISbox_in05_9770, s_out => Sout09_9848, clk => clk, reset => reset); 
    -- logger for split-operator call_stmt_9851_call flow-through 
    process(Sout14_9851) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:call_stmt_9851_call:flowthrough inputs: " & " ISbox_in06_9776 = "& Convert_SLV_To_Hex_String(ISbox_in06_9776) & " outputs:" & " Sout14_9851= "  & Convert_SLV_To_Hex_String(Sout14_9851));
      --
    end process; 
    call_inst_11896: Inv_Sbox_3_Volatile port map(s_in => ISbox_in06_9776, s_out => Sout14_9851, clk => clk, reset => reset); 
    -- logger for split-operator call_stmt_9854_call flow-through 
    process(Sout03_9854) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:call_stmt_9854_call:flowthrough inputs: " & " ISbox_in07_9782 = "& Convert_SLV_To_Hex_String(ISbox_in07_9782) & " outputs:" & " Sout03_9854= "  & Convert_SLV_To_Hex_String(Sout03_9854));
      --
    end process; 
    call_inst_11897: Inv_Sbox_4_Volatile port map(s_in => ISbox_in07_9782, s_out => Sout03_9854, clk => clk, reset => reset); 
    -- logger for split-operator call_stmt_9857_call flow-through 
    process(Sout08_9857) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:call_stmt_9857_call:flowthrough inputs: " & " ISbox_in08_9788 = "& Convert_SLV_To_Hex_String(ISbox_in08_9788) & " outputs:" & " Sout08_9857= "  & Convert_SLV_To_Hex_String(Sout08_9857));
      --
    end process; 
    call_inst_11898: Inv_Sbox_1_Volatile port map(s_in => ISbox_in08_9788, s_out => Sout08_9857, clk => clk, reset => reset); 
    -- logger for split-operator call_stmt_9860_call flow-through 
    process(Sout13_9860) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:call_stmt_9860_call:flowthrough inputs: " & " ISbox_in09_9794 = "& Convert_SLV_To_Hex_String(ISbox_in09_9794) & " outputs:" & " Sout13_9860= "  & Convert_SLV_To_Hex_String(Sout13_9860));
      --
    end process; 
    call_inst_11899: Inv_Sbox_2_Volatile port map(s_in => ISbox_in09_9794, s_out => Sout13_9860, clk => clk, reset => reset); 
    -- logger for split-operator call_stmt_9863_call flow-through 
    process(Sout02_9863) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:call_stmt_9863_call:flowthrough inputs: " & " ISbox_in10_9800 = "& Convert_SLV_To_Hex_String(ISbox_in10_9800) & " outputs:" & " Sout02_9863= "  & Convert_SLV_To_Hex_String(Sout02_9863));
      --
    end process; 
    call_inst_11900: Inv_Sbox_3_Volatile port map(s_in => ISbox_in10_9800, s_out => Sout02_9863, clk => clk, reset => reset); 
    -- logger for split-operator call_stmt_9866_call flow-through 
    process(Sout07_9866) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:call_stmt_9866_call:flowthrough inputs: " & " ISbox_in11_9806 = "& Convert_SLV_To_Hex_String(ISbox_in11_9806) & " outputs:" & " Sout07_9866= "  & Convert_SLV_To_Hex_String(Sout07_9866));
      --
    end process; 
    call_inst_11901: Inv_Sbox_4_Volatile port map(s_in => ISbox_in11_9806, s_out => Sout07_9866, clk => clk, reset => reset); 
    -- logger for split-operator call_stmt_9869_call flow-through 
    process(Sout12_9869) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:call_stmt_9869_call:flowthrough inputs: " & " ISbox_in12_9812 = "& Convert_SLV_To_Hex_String(ISbox_in12_9812) & " outputs:" & " Sout12_9869= "  & Convert_SLV_To_Hex_String(Sout12_9869));
      --
    end process; 
    call_inst_11902: Inv_Sbox_1_Volatile port map(s_in => ISbox_in12_9812, s_out => Sout12_9869, clk => clk, reset => reset); 
    -- logger for split-operator call_stmt_9872_call flow-through 
    process(Sout01_9872) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:call_stmt_9872_call:flowthrough inputs: " & " ISbox_in13_9818 = "& Convert_SLV_To_Hex_String(ISbox_in13_9818) & " outputs:" & " Sout01_9872= "  & Convert_SLV_To_Hex_String(Sout01_9872));
      --
    end process; 
    call_inst_11903: Inv_Sbox_2_Volatile port map(s_in => ISbox_in13_9818, s_out => Sout01_9872, clk => clk, reset => reset); 
    -- logger for split-operator call_stmt_9875_call flow-through 
    process(Sout06_9875) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:call_stmt_9875_call:flowthrough inputs: " & " ISbox_in14_9824 = "& Convert_SLV_To_Hex_String(ISbox_in14_9824) & " outputs:" & " Sout06_9875= "  & Convert_SLV_To_Hex_String(Sout06_9875));
      --
    end process; 
    call_inst_11904: Inv_Sbox_3_Volatile port map(s_in => ISbox_in14_9824, s_out => Sout06_9875, clk => clk, reset => reset); 
    -- logger for split-operator call_stmt_9878_call flow-through 
    process(Sout11_9878) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:dec_round:DP:call_stmt_9878_call:flowthrough inputs: " & " ISbox_in15_9830 = "& Convert_SLV_To_Hex_String(ISbox_in15_9830) & " outputs:" & " Sout11_9878= "  & Convert_SLV_To_Hex_String(Sout11_9878));
      --
    end process; 
    call_inst_11905: Inv_Sbox_4_Volatile port map(s_in => ISbox_in15_9830, s_out => Sout11_9878, clk => clk, reset => reset); 
    -- 
  end Block; -- data_path
  -- 
end dec_round_Operator_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library GhdlLink;
use GhdlLink.LogUtilities.all;
library work;
use work.ahir_system_global_package.all;
entity ahir_system is  -- system 
  port (-- 
    clk : in std_logic;
    reset : in std_logic;
    in_data_pipe_write_data: in std_logic_vector(63 downto 0);
    in_data_pipe_write_req : in std_logic_vector(0 downto 0);
    in_data_pipe_write_ack : out std_logic_vector(0 downto 0);
    out_data_pipe_read_data: out std_logic_vector(63 downto 0);
    out_data_pipe_read_req : in std_logic_vector(0 downto 0);
    out_data_pipe_read_ack : out std_logic_vector(0 downto 0)); -- 
  -- 
end entity; 
architecture ahir_system_arch  of ahir_system is -- system-architecture 
  -- declarations related to module Inv_Sbox_1
  -- declarations related to module Inv_Sbox_2
  -- declarations related to module Inv_Sbox_3
  -- declarations related to module Inv_Sbox_4
  -- declarations related to module MUL2
  -- declarations related to module c_block_daemon_in
  component c_block_daemon_in is -- 
    generic (tag_length : integer); 
    port ( -- 
      in_data_pipe_read_req : out  std_logic_vector(0 downto 0);
      in_data_pipe_read_ack : in   std_logic_vector(0 downto 0);
      in_data_pipe_read_data : in   std_logic_vector(63 downto 0);
      in_buf_pipe_write_req : out  std_logic_vector(0 downto 0);
      in_buf_pipe_write_ack : in   std_logic_vector(0 downto 0);
      in_buf_pipe_write_data : out  std_logic_vector(127 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module c_block_daemon_in
  signal c_block_daemon_in_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal c_block_daemon_in_tag_out   : std_logic_vector(1 downto 0);
  signal c_block_daemon_in_start_req : std_logic;
  signal c_block_daemon_in_start_ack : std_logic;
  signal c_block_daemon_in_fin_req   : std_logic;
  signal c_block_daemon_in_fin_ack : std_logic;
  -- declarations related to module c_block_daemon_out
  component c_block_daemon_out is -- 
    generic (tag_length : integer); 
    port ( -- 
      out_buf_pipe_read_req : out  std_logic_vector(0 downto 0);
      out_buf_pipe_read_ack : in   std_logic_vector(0 downto 0);
      out_buf_pipe_read_data : in   std_logic_vector(127 downto 0);
      out_data_pipe_write_req : out  std_logic_vector(0 downto 0);
      out_data_pipe_write_ack : in   std_logic_vector(0 downto 0);
      out_data_pipe_write_data : out  std_logic_vector(63 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module c_block_daemon_out
  signal c_block_daemon_out_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal c_block_daemon_out_tag_out   : std_logic_vector(1 downto 0);
  signal c_block_daemon_out_start_req : std_logic;
  signal c_block_daemon_out_start_ack : std_logic;
  signal c_block_daemon_out_fin_req   : std_logic;
  signal c_block_daemon_out_fin_ack : std_logic;
  -- declarations related to module d_block_daemon
  component d_block_daemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      in_buf_pipe_read_req : out  std_logic_vector(0 downto 0);
      in_buf_pipe_read_ack : in   std_logic_vector(0 downto 0);
      in_buf_pipe_read_data : in   std_logic_vector(127 downto 0);
      out_buf_pipe_write_req : out  std_logic_vector(0 downto 0);
      out_buf_pipe_write_ack : in   std_logic_vector(0 downto 0);
      out_buf_pipe_write_data : out  std_logic_vector(127 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module d_block_daemon
  signal d_block_daemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal d_block_daemon_tag_out   : std_logic_vector(1 downto 0);
  signal d_block_daemon_start_req : std_logic;
  signal d_block_daemon_start_ack : std_logic;
  signal d_block_daemon_fin_req   : std_logic;
  signal d_block_daemon_fin_ack : std_logic;
  -- declarations related to module dec_round
  -- aggregate signals for write to pipe in_buf
  signal in_buf_pipe_write_data: std_logic_vector(127 downto 0);
  signal in_buf_pipe_write_req: std_logic_vector(0 downto 0);
  signal in_buf_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe in_buf
  signal in_buf_pipe_read_data: std_logic_vector(127 downto 0);
  signal in_buf_pipe_read_req: std_logic_vector(0 downto 0);
  signal in_buf_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe in_data
  signal in_data_pipe_read_data: std_logic_vector(63 downto 0);
  signal in_data_pipe_read_req: std_logic_vector(0 downto 0);
  signal in_data_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe out_buf
  signal out_buf_pipe_write_data: std_logic_vector(127 downto 0);
  signal out_buf_pipe_write_req: std_logic_vector(0 downto 0);
  signal out_buf_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe out_buf
  signal out_buf_pipe_read_data: std_logic_vector(127 downto 0);
  signal out_buf_pipe_read_req: std_logic_vector(0 downto 0);
  signal out_buf_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe out_data
  signal out_data_pipe_write_data: std_logic_vector(63 downto 0);
  signal out_data_pipe_write_req: std_logic_vector(0 downto 0);
  signal out_data_pipe_write_ack: std_logic_vector(0 downto 0);
  -- 
begin -- 
  -- module c_block_daemon_in
  c_block_daemon_in_instance:c_block_daemon_in-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => c_block_daemon_in_start_req,
      start_ack => c_block_daemon_in_start_ack,
      fin_req => c_block_daemon_in_fin_req,
      fin_ack => c_block_daemon_in_fin_ack,
      clk => clk,
      reset => reset,
      in_data_pipe_read_req => in_data_pipe_read_req(0 downto 0),
      in_data_pipe_read_ack => in_data_pipe_read_ack(0 downto 0),
      in_data_pipe_read_data => in_data_pipe_read_data(63 downto 0),
      in_buf_pipe_write_req => in_buf_pipe_write_req(0 downto 0),
      in_buf_pipe_write_ack => in_buf_pipe_write_ack(0 downto 0),
      in_buf_pipe_write_data => in_buf_pipe_write_data(127 downto 0),
      tag_in => c_block_daemon_in_tag_in,
      tag_out => c_block_daemon_in_tag_out-- 
    ); -- 
  -- module will be run forever 
  c_block_daemon_in_tag_in <= (others => '0');
  c_block_daemon_in_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => c_block_daemon_in_start_req, start_ack => c_block_daemon_in_start_ack,  fin_req => c_block_daemon_in_fin_req,  fin_ack => c_block_daemon_in_fin_ack);
  -- module c_block_daemon_out
  c_block_daemon_out_instance:c_block_daemon_out-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => c_block_daemon_out_start_req,
      start_ack => c_block_daemon_out_start_ack,
      fin_req => c_block_daemon_out_fin_req,
      fin_ack => c_block_daemon_out_fin_ack,
      clk => clk,
      reset => reset,
      out_buf_pipe_read_req => out_buf_pipe_read_req(0 downto 0),
      out_buf_pipe_read_ack => out_buf_pipe_read_ack(0 downto 0),
      out_buf_pipe_read_data => out_buf_pipe_read_data(127 downto 0),
      out_data_pipe_write_req => out_data_pipe_write_req(0 downto 0),
      out_data_pipe_write_ack => out_data_pipe_write_ack(0 downto 0),
      out_data_pipe_write_data => out_data_pipe_write_data(63 downto 0),
      tag_in => c_block_daemon_out_tag_in,
      tag_out => c_block_daemon_out_tag_out-- 
    ); -- 
  -- module will be run forever 
  c_block_daemon_out_tag_in <= (others => '0');
  c_block_daemon_out_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => c_block_daemon_out_start_req, start_ack => c_block_daemon_out_start_ack,  fin_req => c_block_daemon_out_fin_req,  fin_ack => c_block_daemon_out_fin_ack);
  -- module d_block_daemon
  d_block_daemon_instance:d_block_daemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => d_block_daemon_start_req,
      start_ack => d_block_daemon_start_ack,
      fin_req => d_block_daemon_fin_req,
      fin_ack => d_block_daemon_fin_ack,
      clk => clk,
      reset => reset,
      in_buf_pipe_read_req => in_buf_pipe_read_req(0 downto 0),
      in_buf_pipe_read_ack => in_buf_pipe_read_ack(0 downto 0),
      in_buf_pipe_read_data => in_buf_pipe_read_data(127 downto 0),
      out_buf_pipe_write_req => out_buf_pipe_write_req(0 downto 0),
      out_buf_pipe_write_ack => out_buf_pipe_write_ack(0 downto 0),
      out_buf_pipe_write_data => out_buf_pipe_write_data(127 downto 0),
      tag_in => d_block_daemon_tag_in,
      tag_out => d_block_daemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  d_block_daemon_tag_in <= (others => '0');
  d_block_daemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => d_block_daemon_start_req, start_ack => d_block_daemon_start_ack,  fin_req => d_block_daemon_fin_req,  fin_ack => d_block_daemon_fin_ack);
  in_buf_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe in_buf",
      num_reads => 1,
      num_writes => 1,
      data_width => 128,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      depth => 256 --
    )
    port map( -- 
      read_req => in_buf_pipe_read_req,
      read_ack => in_buf_pipe_read_ack,
      read_data => in_buf_pipe_read_data,
      write_req => in_buf_pipe_write_req,
      write_ack => in_buf_pipe_write_ack,
      write_data => in_buf_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  in_data_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe in_data",
      num_reads => 1,
      num_writes => 1,
      data_width => 64,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      depth => 2 --
    )
    port map( -- 
      read_req => in_data_pipe_read_req,
      read_ack => in_data_pipe_read_ack,
      read_data => in_data_pipe_read_data,
      write_req => in_data_pipe_write_req,
      write_ack => in_data_pipe_write_ack,
      write_data => in_data_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  out_buf_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe out_buf",
      num_reads => 1,
      num_writes => 1,
      data_width => 128,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      depth => 256 --
    )
    port map( -- 
      read_req => out_buf_pipe_read_req,
      read_ack => out_buf_pipe_read_ack,
      read_data => out_buf_pipe_read_data,
      write_req => out_buf_pipe_write_req,
      write_ack => out_buf_pipe_write_ack,
      write_data => out_buf_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  out_data_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe out_data",
      num_reads => 1,
      num_writes => 1,
      data_width => 64,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      depth => 2 --
    )
    port map( -- 
      read_req => out_data_pipe_read_req,
      read_ack => out_data_pipe_read_ack,
      read_data => out_data_pipe_read_data,
      write_req => out_data_pipe_write_req,
      write_ack => out_data_pipe_write_ack,
      write_data => out_data_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- 
end ahir_system_arch;
