-- VHDL produced by vc2vhdl from virtual circuit (vc) description 
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library work;
use work.ahir_system_global_package.all;
entity In_wrap_daemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    w_in_buf_pipe_read_req : out  std_logic_vector(0 downto 0);
    w_in_buf_pipe_read_ack : in   std_logic_vector(0 downto 0);
    w_in_buf_pipe_read_data : in   std_logic_vector(127 downto 0);
    cmd_in_pipe_write_req : out  std_logic_vector(0 downto 0);
    cmd_in_pipe_write_ack : in   std_logic_vector(0 downto 0);
    cmd_in_pipe_write_data : out  std_logic_vector(63 downto 0);
    d_in_buf_pipe_write_req : out  std_logic_vector(0 downto 0);
    d_in_buf_pipe_write_ack : in   std_logic_vector(0 downto 0);
    d_in_buf_pipe_write_data : out  std_logic_vector(127 downto 0);
    e_in_buf_pipe_write_req : out  std_logic_vector(0 downto 0);
    e_in_buf_pipe_write_ack : in   std_logic_vector(0 downto 0);
    e_in_buf_pipe_write_data : out  std_logic_vector(127 downto 0);
    out_wrap_cmd_pipe_write_req : out  std_logic_vector(0 downto 0);
    out_wrap_cmd_pipe_write_ack : in   std_logic_vector(0 downto 0);
    out_wrap_cmd_pipe_write_data : out  std_logic_vector(63 downto 0);
    out_wrap_data_pipe_write_req : out  std_logic_vector(0 downto 0);
    out_wrap_data_pipe_write_ack : in   std_logic_vector(0 downto 0);
    out_wrap_data_pipe_write_data : out  std_logic_vector(127 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity In_wrap_daemon;
architecture In_wrap_daemon_arch of In_wrap_daemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal In_wrap_daemon_CP_0_start: Boolean;
  signal In_wrap_daemon_CP_0_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal RPIPE_w_in_buf_33_inst_req_0 : boolean;
  signal RPIPE_w_in_buf_33_inst_ack_0 : boolean;
  signal RPIPE_w_in_buf_33_inst_req_1 : boolean;
  signal RPIPE_w_in_buf_33_inst_ack_1 : boolean;
  signal WPIPE_cmd_in_43_inst_req_0 : boolean;
  signal WPIPE_cmd_in_43_inst_ack_0 : boolean;
  signal WPIPE_cmd_in_43_inst_req_1 : boolean;
  signal WPIPE_cmd_in_43_inst_ack_1 : boolean;
  signal WPIPE_out_wrap_cmd_46_inst_req_0 : boolean;
  signal WPIPE_out_wrap_cmd_46_inst_ack_0 : boolean;
  signal WPIPE_out_wrap_cmd_46_inst_req_1 : boolean;
  signal WPIPE_out_wrap_cmd_46_inst_ack_1 : boolean;
  signal WPIPE_cmd_in_89_inst_req_0 : boolean;
  signal WPIPE_cmd_in_89_inst_ack_0 : boolean;
  signal WPIPE_cmd_in_89_inst_req_1 : boolean;
  signal WPIPE_cmd_in_89_inst_ack_1 : boolean;
  signal if_stmt_71_branch_req_0 : boolean;
  signal if_stmt_71_branch_ack_1 : boolean;
  signal if_stmt_71_branch_ack_0 : boolean;
  signal RPIPE_w_in_buf_76_inst_req_0 : boolean;
  signal RPIPE_w_in_buf_76_inst_ack_0 : boolean;
  signal RPIPE_w_in_buf_76_inst_req_1 : boolean;
  signal RPIPE_w_in_buf_76_inst_ack_1 : boolean;
  signal slice_80_inst_req_0 : boolean;
  signal slice_80_inst_ack_0 : boolean;
  signal slice_80_inst_req_1 : boolean;
  signal slice_80_inst_ack_1 : boolean;
  signal slice_84_inst_req_0 : boolean;
  signal slice_84_inst_ack_0 : boolean;
  signal slice_84_inst_req_1 : boolean;
  signal slice_84_inst_ack_1 : boolean;
  signal WPIPE_cmd_in_86_inst_req_0 : boolean;
  signal WPIPE_cmd_in_86_inst_ack_0 : boolean;
  signal WPIPE_cmd_in_86_inst_req_1 : boolean;
  signal WPIPE_cmd_in_86_inst_ack_1 : boolean;
  signal n_count_var2_154_145_buf_req_1 : boolean;
  signal n_count_var2_154_145_buf_ack_1 : boolean;
  signal phi_stmt_142_req_1 : boolean;
  signal phi_stmt_142_ack_0 : boolean;
  signal phi_stmt_109_req_0 : boolean;
  signal OR_u15_u15_106_inst_req_0 : boolean;
  signal OR_u15_u15_106_inst_ack_0 : boolean;
  signal OR_u15_u15_106_inst_req_1 : boolean;
  signal OR_u15_u15_106_inst_ack_1 : boolean;
  signal if_stmt_114_branch_req_0 : boolean;
  signal if_stmt_114_branch_ack_1 : boolean;
  signal if_stmt_114_branch_ack_0 : boolean;
  signal RPIPE_w_in_buf_119_inst_req_0 : boolean;
  signal RPIPE_w_in_buf_119_inst_ack_0 : boolean;
  signal RPIPE_w_in_buf_119_inst_req_1 : boolean;
  signal RPIPE_w_in_buf_119_inst_ack_1 : boolean;
  signal WPIPE_e_in_buf_118_inst_req_0 : boolean;
  signal WPIPE_e_in_buf_118_inst_ack_0 : boolean;
  signal WPIPE_e_in_buf_118_inst_req_1 : boolean;
  signal WPIPE_e_in_buf_118_inst_ack_1 : boolean;
  signal RPIPE_w_in_buf_123_inst_req_0 : boolean;
  signal RPIPE_w_in_buf_123_inst_ack_0 : boolean;
  signal RPIPE_w_in_buf_123_inst_req_1 : boolean;
  signal RPIPE_w_in_buf_123_inst_ack_1 : boolean;
  signal WPIPE_d_in_buf_122_inst_req_0 : boolean;
  signal WPIPE_d_in_buf_122_inst_ack_0 : boolean;
  signal WPIPE_d_in_buf_122_inst_req_1 : boolean;
  signal WPIPE_d_in_buf_122_inst_ack_1 : boolean;
  signal if_stmt_131_branch_req_0 : boolean;
  signal if_stmt_131_branch_ack_1 : boolean;
  signal if_stmt_131_branch_ack_0 : boolean;
  signal if_stmt_137_branch_req_0 : boolean;
  signal if_stmt_137_branch_ack_1 : boolean;
  signal if_stmt_137_branch_ack_0 : boolean;
  signal RPIPE_w_in_buf_148_inst_req_0 : boolean;
  signal RPIPE_w_in_buf_148_inst_ack_0 : boolean;
  signal RPIPE_w_in_buf_148_inst_req_1 : boolean;
  signal RPIPE_w_in_buf_148_inst_ack_1 : boolean;
  signal WPIPE_out_wrap_data_147_inst_req_0 : boolean;
  signal WPIPE_out_wrap_data_147_inst_ack_0 : boolean;
  signal WPIPE_out_wrap_data_147_inst_req_1 : boolean;
  signal WPIPE_out_wrap_data_147_inst_ack_1 : boolean;
  signal if_stmt_155_branch_req_0 : boolean;
  signal if_stmt_155_branch_ack_1 : boolean;
  signal if_stmt_155_branch_ack_0 : boolean;
  signal n_count_var_130_144_buf_req_0 : boolean;
  signal n_count_var_130_144_buf_ack_0 : boolean;
  signal n_count_var_130_144_buf_req_1 : boolean;
  signal n_count_var_130_144_buf_ack_1 : boolean;
  signal phi_stmt_142_req_0 : boolean;
  signal n_count_var2_154_145_buf_req_0 : boolean;
  signal n_count_var2_154_145_buf_ack_0 : boolean;
  signal n_count_var_130_112_buf_req_0 : boolean;
  signal n_count_var_130_112_buf_ack_0 : boolean;
  signal n_count_var_130_112_buf_req_1 : boolean;
  signal n_count_var_130_112_buf_ack_1 : boolean;
  signal phi_stmt_109_req_1 : boolean;
  signal phi_stmt_109_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "In_wrap_daemon_input_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      bypass_flag => true,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  In_wrap_daemon_CP_0_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "In_wrap_daemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= In_wrap_daemon_CP_0_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= In_wrap_daemon_CP_0_start & tag_ilock_write_ack_symbol;
    gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= In_wrap_daemon_CP_0_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  In_wrap_daemon_CP_0: Block -- control-path 
    signal In_wrap_daemon_CP_0_elements: BooleanArray(132 downto 0);
    -- 
  begin -- 
    In_wrap_daemon_CP_0_elements(0) <= In_wrap_daemon_CP_0_start;
    In_wrap_daemon_CP_0_symbol <= In_wrap_daemon_CP_0_elements(132);
    -- CP-element group 0:  transition  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (2) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_31/$entry
      -- 
    -- CP-element group 1:  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	12 
    -- CP-element group 1:  members (2) 
      -- CP-element group 1: 	 branch_block_stmt_31/branch_block_stmt_31__entry__
      -- CP-element group 1: 	 branch_block_stmt_31/assign_stmt_34__entry__
      -- 
    In_wrap_daemon_CP_0_elements(1) <= In_wrap_daemon_CP_0_elements(0);
    -- CP-element group 2:  place  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	14 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	15 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_31/assign_stmt_34__exit__
      -- CP-element group 2: 	 branch_block_stmt_31/assign_stmt_38_to_assign_stmt_42__entry__
      -- 
    In_wrap_daemon_CP_0_elements(2) <= In_wrap_daemon_CP_0_elements(14);
    -- CP-element group 3:  place  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	15 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	16 
    -- CP-element group 3:  members (2) 
      -- CP-element group 3: 	 branch_block_stmt_31/assign_stmt_38_to_assign_stmt_42__exit__
      -- CP-element group 3: 	 branch_block_stmt_31/assign_stmt_45__entry__
      -- 
    In_wrap_daemon_CP_0_elements(3) <= In_wrap_daemon_CP_0_elements(15);
    -- CP-element group 4:  place  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	18 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	19 
    -- CP-element group 4:  members (2) 
      -- CP-element group 4: 	 branch_block_stmt_31/assign_stmt_45__exit__
      -- CP-element group 4: 	 branch_block_stmt_31/assign_stmt_48__entry__
      -- 
    In_wrap_daemon_CP_0_elements(4) <= In_wrap_daemon_CP_0_elements(18);
    -- CP-element group 5:  place  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	21 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	22 
    -- CP-element group 5:  members (2) 
      -- CP-element group 5: 	 branch_block_stmt_31/assign_stmt_48__exit__
      -- CP-element group 5: 	 branch_block_stmt_31/assign_stmt_52_to_assign_stmt_70__entry__
      -- 
    In_wrap_daemon_CP_0_elements(5) <= In_wrap_daemon_CP_0_elements(21);
    -- CP-element group 6:  branch  place  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	22 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	23 
    -- CP-element group 6: 	24 
    -- CP-element group 6:  members (2) 
      -- CP-element group 6: 	 branch_block_stmt_31/assign_stmt_52_to_assign_stmt_70__exit__
      -- CP-element group 6: 	 branch_block_stmt_31/if_stmt_71__entry__
      -- 
    In_wrap_daemon_CP_0_elements(6) <= In_wrap_daemon_CP_0_elements(22);
    -- CP-element group 7:  merge  place  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	29 
    -- CP-element group 7: 	34 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	50 
    -- CP-element group 7:  members (2) 
      -- CP-element group 7: 	 branch_block_stmt_31/if_stmt_71__exit__
      -- CP-element group 7: 	 branch_block_stmt_31/assign_stmt_107__entry__
      -- 
    In_wrap_daemon_CP_0_elements(7) <= OrReduce(In_wrap_daemon_CP_0_elements(29) & In_wrap_daemon_CP_0_elements(34));
    -- CP-element group 8:  branch  place  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	52 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	123 
    -- CP-element group 8: 	124 
    -- CP-element group 8:  members (2) 
      -- CP-element group 8: 	 branch_block_stmt_31/assign_stmt_107__exit__
      -- CP-element group 8: 	 branch_block_stmt_31/merge_stmt_108__entry__
      -- 
    In_wrap_daemon_CP_0_elements(8) <= In_wrap_daemon_CP_0_elements(52);
    -- CP-element group 9:  merge  branch  place  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	131 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	53 
    -- CP-element group 9: 	54 
    -- CP-element group 9:  members (2) 
      -- CP-element group 9: 	 branch_block_stmt_31/merge_stmt_108__exit__
      -- CP-element group 9: 	 branch_block_stmt_31/if_stmt_114__entry__
      -- 
    In_wrap_daemon_CP_0_elements(9) <= In_wrap_daemon_CP_0_elements(131);
    -- CP-element group 10:  merge  place  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	61 
    -- CP-element group 10: 	68 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	74 
    -- CP-element group 10:  members (2) 
      -- CP-element group 10: 	 branch_block_stmt_31/if_stmt_114__exit__
      -- CP-element group 10: 	 branch_block_stmt_31/assign_stmt_130__entry__
      -- 
    In_wrap_daemon_CP_0_elements(10) <= OrReduce(In_wrap_daemon_CP_0_elements(61) & In_wrap_daemon_CP_0_elements(68));
    -- CP-element group 11:  branch  place  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	74 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	75 
    -- CP-element group 11: 	76 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_31/assign_stmt_130__exit__
      -- CP-element group 11: 	 branch_block_stmt_31/if_stmt_131__entry__
      -- 
    In_wrap_daemon_CP_0_elements(11) <= In_wrap_daemon_CP_0_elements(74);
    -- CP-element group 12:  transition  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	1 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (4) 
      -- CP-element group 12: 	 branch_block_stmt_31/assign_stmt_34/RPIPE_w_in_buf_33_Sample/$entry
      -- CP-element group 12: 	 branch_block_stmt_31/assign_stmt_34/$entry
      -- CP-element group 12: 	 branch_block_stmt_31/assign_stmt_34/RPIPE_w_in_buf_33_sample_start_
      -- CP-element group 12: 	 branch_block_stmt_31/assign_stmt_34/RPIPE_w_in_buf_33_Sample/rr
      -- 
    rr_40_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_40_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => In_wrap_daemon_CP_0_elements(12), ack => RPIPE_w_in_buf_33_inst_req_0); -- 
    In_wrap_daemon_CP_0_elements(12) <= In_wrap_daemon_CP_0_elements(1);
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_31/assign_stmt_34/RPIPE_w_in_buf_33_Sample/$exit
      -- CP-element group 13: 	 branch_block_stmt_31/assign_stmt_34/RPIPE_w_in_buf_33_sample_completed_
      -- CP-element group 13: 	 branch_block_stmt_31/assign_stmt_34/RPIPE_w_in_buf_33_update_start_
      -- CP-element group 13: 	 branch_block_stmt_31/assign_stmt_34/RPIPE_w_in_buf_33_Sample/ra
      -- CP-element group 13: 	 branch_block_stmt_31/assign_stmt_34/RPIPE_w_in_buf_33_Update/$entry
      -- CP-element group 13: 	 branch_block_stmt_31/assign_stmt_34/RPIPE_w_in_buf_33_Update/cr
      -- 
    ra_41_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_w_in_buf_33_inst_ack_0, ack => In_wrap_daemon_CP_0_elements(13)); -- 
    cr_45_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_45_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => In_wrap_daemon_CP_0_elements(13), ack => RPIPE_w_in_buf_33_inst_req_1); -- 
    -- CP-element group 14:  transition  input  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	2 
    -- CP-element group 14:  members (4) 
      -- CP-element group 14: 	 branch_block_stmt_31/assign_stmt_34/$exit
      -- CP-element group 14: 	 branch_block_stmt_31/assign_stmt_34/RPIPE_w_in_buf_33_update_completed_
      -- CP-element group 14: 	 branch_block_stmt_31/assign_stmt_34/RPIPE_w_in_buf_33_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_31/assign_stmt_34/RPIPE_w_in_buf_33_Update/ca
      -- 
    ca_46_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_w_in_buf_33_inst_ack_1, ack => In_wrap_daemon_CP_0_elements(14)); -- 
    -- CP-element group 15:  join  fork  transition  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	2 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	3 
    -- CP-element group 15:  members (34) 
      -- CP-element group 15: 	 branch_block_stmt_31/assign_stmt_38_to_assign_stmt_42/$entry
      -- CP-element group 15: 	 branch_block_stmt_31/assign_stmt_38_to_assign_stmt_42/$exit
      -- CP-element group 15: 	 branch_block_stmt_31/assign_stmt_38_to_assign_stmt_42/slice_37_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_31/assign_stmt_38_to_assign_stmt_42/slice_37_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_31/assign_stmt_38_to_assign_stmt_42/slice_37_update_start_
      -- CP-element group 15: 	 branch_block_stmt_31/assign_stmt_38_to_assign_stmt_42/slice_37_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_31/assign_stmt_38_to_assign_stmt_42/R_head_in_36_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_31/assign_stmt_38_to_assign_stmt_42/R_head_in_36_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_31/assign_stmt_38_to_assign_stmt_42/R_head_in_36_update_start_
      -- CP-element group 15: 	 branch_block_stmt_31/assign_stmt_38_to_assign_stmt_42/R_head_in_36_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_31/assign_stmt_38_to_assign_stmt_42/slice_41_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_31/assign_stmt_38_to_assign_stmt_42/slice_41_Update/ca
      -- CP-element group 15: 	 branch_block_stmt_31/assign_stmt_38_to_assign_stmt_42/slice_37_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_31/assign_stmt_38_to_assign_stmt_42/slice_37_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_31/assign_stmt_38_to_assign_stmt_42/slice_37_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_31/assign_stmt_38_to_assign_stmt_42/slice_37_Sample/ra
      -- CP-element group 15: 	 branch_block_stmt_31/assign_stmt_38_to_assign_stmt_42/slice_37_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_31/assign_stmt_38_to_assign_stmt_42/slice_37_Update/$exit
      -- CP-element group 15: 	 branch_block_stmt_31/assign_stmt_38_to_assign_stmt_42/slice_37_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_31/assign_stmt_38_to_assign_stmt_42/slice_37_Update/ca
      -- CP-element group 15: 	 branch_block_stmt_31/assign_stmt_38_to_assign_stmt_42/slice_41_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_31/assign_stmt_38_to_assign_stmt_42/slice_41_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_31/assign_stmt_38_to_assign_stmt_42/slice_41_update_start_
      -- CP-element group 15: 	 branch_block_stmt_31/assign_stmt_38_to_assign_stmt_42/slice_41_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_31/assign_stmt_38_to_assign_stmt_42/R_head_in_40_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_31/assign_stmt_38_to_assign_stmt_42/R_head_in_40_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_31/assign_stmt_38_to_assign_stmt_42/R_head_in_40_update_start_
      -- CP-element group 15: 	 branch_block_stmt_31/assign_stmt_38_to_assign_stmt_42/R_head_in_40_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_31/assign_stmt_38_to_assign_stmt_42/slice_41_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_31/assign_stmt_38_to_assign_stmt_42/slice_41_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_31/assign_stmt_38_to_assign_stmt_42/slice_41_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_31/assign_stmt_38_to_assign_stmt_42/slice_41_Sample/ra
      -- CP-element group 15: 	 branch_block_stmt_31/assign_stmt_38_to_assign_stmt_42/slice_41_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_31/assign_stmt_38_to_assign_stmt_42/slice_41_Update/$exit
      -- 
    In_wrap_daemon_CP_0_elements(15) <= In_wrap_daemon_CP_0_elements(2);
    -- CP-element group 16:  transition  output  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	3 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	17 
    -- CP-element group 16:  members (8) 
      -- CP-element group 16: 	 branch_block_stmt_31/assign_stmt_45/$entry
      -- CP-element group 16: 	 branch_block_stmt_31/assign_stmt_45/R_head1_44_sample_start_
      -- CP-element group 16: 	 branch_block_stmt_31/assign_stmt_45/R_head1_44_sample_completed_
      -- CP-element group 16: 	 branch_block_stmt_31/assign_stmt_45/R_head1_44_update_start_
      -- CP-element group 16: 	 branch_block_stmt_31/assign_stmt_45/R_head1_44_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_31/assign_stmt_45/WPIPE_cmd_in_43_sample_start_
      -- CP-element group 16: 	 branch_block_stmt_31/assign_stmt_45/WPIPE_cmd_in_43_Sample/$entry
      -- CP-element group 16: 	 branch_block_stmt_31/assign_stmt_45/WPIPE_cmd_in_43_Sample/req
      -- 
    req_100_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_100_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => In_wrap_daemon_CP_0_elements(16), ack => WPIPE_cmd_in_43_inst_req_0); -- 
    In_wrap_daemon_CP_0_elements(16) <= In_wrap_daemon_CP_0_elements(3);
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	16 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_31/assign_stmt_45/WPIPE_cmd_in_43_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_31/assign_stmt_45/WPIPE_cmd_in_43_update_start_
      -- CP-element group 17: 	 branch_block_stmt_31/assign_stmt_45/WPIPE_cmd_in_43_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_31/assign_stmt_45/WPIPE_cmd_in_43_Sample/ack
      -- CP-element group 17: 	 branch_block_stmt_31/assign_stmt_45/WPIPE_cmd_in_43_Update/$entry
      -- CP-element group 17: 	 branch_block_stmt_31/assign_stmt_45/WPIPE_cmd_in_43_Update/req
      -- 
    ack_101_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_cmd_in_43_inst_ack_0, ack => In_wrap_daemon_CP_0_elements(17)); -- 
    req_105_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_105_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => In_wrap_daemon_CP_0_elements(17), ack => WPIPE_cmd_in_43_inst_req_1); -- 
    -- CP-element group 18:  transition  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	4 
    -- CP-element group 18:  members (4) 
      -- CP-element group 18: 	 branch_block_stmt_31/assign_stmt_45/$exit
      -- CP-element group 18: 	 branch_block_stmt_31/assign_stmt_45/WPIPE_cmd_in_43_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_31/assign_stmt_45/WPIPE_cmd_in_43_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_31/assign_stmt_45/WPIPE_cmd_in_43_Update/ack
      -- 
    ack_106_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_cmd_in_43_inst_ack_1, ack => In_wrap_daemon_CP_0_elements(18)); -- 
    -- CP-element group 19:  transition  output  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	4 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19:  members (8) 
      -- CP-element group 19: 	 branch_block_stmt_31/assign_stmt_48/$entry
      -- CP-element group 19: 	 branch_block_stmt_31/assign_stmt_48/R_head1_47_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_31/assign_stmt_48/R_head1_47_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_31/assign_stmt_48/R_head1_47_update_start_
      -- CP-element group 19: 	 branch_block_stmt_31/assign_stmt_48/R_head1_47_update_completed_
      -- CP-element group 19: 	 branch_block_stmt_31/assign_stmt_48/WPIPE_out_wrap_cmd_46_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_31/assign_stmt_48/WPIPE_out_wrap_cmd_46_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_31/assign_stmt_48/WPIPE_out_wrap_cmd_46_Sample/req
      -- 
    req_121_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_121_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => In_wrap_daemon_CP_0_elements(19), ack => WPIPE_out_wrap_cmd_46_inst_req_0); -- 
    In_wrap_daemon_CP_0_elements(19) <= In_wrap_daemon_CP_0_elements(4);
    -- CP-element group 20:  transition  input  output  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	21 
    -- CP-element group 20:  members (6) 
      -- CP-element group 20: 	 branch_block_stmt_31/assign_stmt_48/WPIPE_out_wrap_cmd_46_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_31/assign_stmt_48/WPIPE_out_wrap_cmd_46_update_start_
      -- CP-element group 20: 	 branch_block_stmt_31/assign_stmt_48/WPIPE_out_wrap_cmd_46_Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_31/assign_stmt_48/WPIPE_out_wrap_cmd_46_Sample/ack
      -- CP-element group 20: 	 branch_block_stmt_31/assign_stmt_48/WPIPE_out_wrap_cmd_46_Update/$entry
      -- CP-element group 20: 	 branch_block_stmt_31/assign_stmt_48/WPIPE_out_wrap_cmd_46_Update/req
      -- 
    ack_122_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_out_wrap_cmd_46_inst_ack_0, ack => In_wrap_daemon_CP_0_elements(20)); -- 
    req_126_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_126_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => In_wrap_daemon_CP_0_elements(20), ack => WPIPE_out_wrap_cmd_46_inst_req_1); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	20 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	5 
    -- CP-element group 21:  members (4) 
      -- CP-element group 21: 	 branch_block_stmt_31/assign_stmt_48/$exit
      -- CP-element group 21: 	 branch_block_stmt_31/assign_stmt_48/WPIPE_out_wrap_cmd_46_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_31/assign_stmt_48/WPIPE_out_wrap_cmd_46_Update/$exit
      -- CP-element group 21: 	 branch_block_stmt_31/assign_stmt_48/WPIPE_out_wrap_cmd_46_Update/ack
      -- 
    ack_127_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_out_wrap_cmd_46_inst_ack_1, ack => In_wrap_daemon_CP_0_elements(21)); -- 
    -- CP-element group 22:  join  fork  transition  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	5 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	6 
    -- CP-element group 22:  members (82) 
      -- CP-element group 22: 	 branch_block_stmt_31/assign_stmt_52_to_assign_stmt_70/slice_60_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_31/assign_stmt_52_to_assign_stmt_70/slice_60_sample_completed_
      -- CP-element group 22: 	 branch_block_stmt_31/assign_stmt_52_to_assign_stmt_70/slice_60_update_start_
      -- CP-element group 22: 	 branch_block_stmt_31/assign_stmt_52_to_assign_stmt_70/$entry
      -- CP-element group 22: 	 branch_block_stmt_31/assign_stmt_52_to_assign_stmt_70/$exit
      -- CP-element group 22: 	 branch_block_stmt_31/assign_stmt_52_to_assign_stmt_70/slice_51_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_31/assign_stmt_52_to_assign_stmt_70/slice_51_sample_completed_
      -- CP-element group 22: 	 branch_block_stmt_31/assign_stmt_52_to_assign_stmt_70/slice_51_update_start_
      -- CP-element group 22: 	 branch_block_stmt_31/assign_stmt_52_to_assign_stmt_70/slice_51_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_31/assign_stmt_52_to_assign_stmt_70/R_head1_50_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_31/assign_stmt_52_to_assign_stmt_70/R_head1_50_sample_completed_
      -- CP-element group 22: 	 branch_block_stmt_31/assign_stmt_52_to_assign_stmt_70/R_head1_50_update_start_
      -- CP-element group 22: 	 branch_block_stmt_31/assign_stmt_52_to_assign_stmt_70/R_head1_50_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_31/assign_stmt_52_to_assign_stmt_70/slice_51_Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_31/assign_stmt_52_to_assign_stmt_70/slice_51_Sample/$exit
      -- CP-element group 22: 	 branch_block_stmt_31/assign_stmt_52_to_assign_stmt_70/slice_51_Sample/rr
      -- CP-element group 22: 	 branch_block_stmt_31/assign_stmt_52_to_assign_stmt_70/slice_51_Sample/ra
      -- CP-element group 22: 	 branch_block_stmt_31/assign_stmt_52_to_assign_stmt_70/slice_51_Update/$entry
      -- CP-element group 22: 	 branch_block_stmt_31/assign_stmt_52_to_assign_stmt_70/slice_51_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_31/assign_stmt_52_to_assign_stmt_70/slice_51_Update/cr
      -- CP-element group 22: 	 branch_block_stmt_31/assign_stmt_52_to_assign_stmt_70/slice_51_Update/ca
      -- CP-element group 22: 	 branch_block_stmt_31/assign_stmt_52_to_assign_stmt_70/slice_56_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_31/assign_stmt_52_to_assign_stmt_70/slice_56_sample_completed_
      -- CP-element group 22: 	 branch_block_stmt_31/assign_stmt_52_to_assign_stmt_70/slice_56_update_start_
      -- CP-element group 22: 	 branch_block_stmt_31/assign_stmt_52_to_assign_stmt_70/slice_56_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_31/assign_stmt_52_to_assign_stmt_70/R_head1_54_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_31/assign_stmt_52_to_assign_stmt_70/R_head1_54_sample_completed_
      -- CP-element group 22: 	 branch_block_stmt_31/assign_stmt_52_to_assign_stmt_70/R_head1_54_update_start_
      -- CP-element group 22: 	 branch_block_stmt_31/assign_stmt_52_to_assign_stmt_70/R_head1_54_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_31/assign_stmt_52_to_assign_stmt_70/slice_56_Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_31/assign_stmt_52_to_assign_stmt_70/slice_56_Sample/$exit
      -- CP-element group 22: 	 branch_block_stmt_31/assign_stmt_52_to_assign_stmt_70/slice_56_Sample/rr
      -- CP-element group 22: 	 branch_block_stmt_31/assign_stmt_52_to_assign_stmt_70/slice_56_Sample/ra
      -- CP-element group 22: 	 branch_block_stmt_31/assign_stmt_52_to_assign_stmt_70/slice_56_Update/$entry
      -- CP-element group 22: 	 branch_block_stmt_31/assign_stmt_52_to_assign_stmt_70/slice_56_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_31/assign_stmt_52_to_assign_stmt_70/slice_56_Update/cr
      -- CP-element group 22: 	 branch_block_stmt_31/assign_stmt_52_to_assign_stmt_70/slice_56_Update/ca
      -- CP-element group 22: 	 branch_block_stmt_31/assign_stmt_52_to_assign_stmt_70/slice_60_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_31/assign_stmt_52_to_assign_stmt_70/R_head1_59_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_31/assign_stmt_52_to_assign_stmt_70/R_head1_59_sample_completed_
      -- CP-element group 22: 	 branch_block_stmt_31/assign_stmt_52_to_assign_stmt_70/R_head1_59_update_start_
      -- CP-element group 22: 	 branch_block_stmt_31/assign_stmt_52_to_assign_stmt_70/R_head1_59_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_31/assign_stmt_52_to_assign_stmt_70/slice_60_Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_31/assign_stmt_52_to_assign_stmt_70/slice_60_Sample/$exit
      -- CP-element group 22: 	 branch_block_stmt_31/assign_stmt_52_to_assign_stmt_70/slice_60_Sample/rr
      -- CP-element group 22: 	 branch_block_stmt_31/assign_stmt_52_to_assign_stmt_70/slice_60_Sample/ra
      -- CP-element group 22: 	 branch_block_stmt_31/assign_stmt_52_to_assign_stmt_70/slice_60_Update/$entry
      -- CP-element group 22: 	 branch_block_stmt_31/assign_stmt_52_to_assign_stmt_70/slice_60_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_31/assign_stmt_52_to_assign_stmt_70/slice_60_Update/cr
      -- CP-element group 22: 	 branch_block_stmt_31/assign_stmt_52_to_assign_stmt_70/slice_60_Update/ca
      -- CP-element group 22: 	 branch_block_stmt_31/assign_stmt_52_to_assign_stmt_70/slice_65_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_31/assign_stmt_52_to_assign_stmt_70/slice_65_sample_completed_
      -- CP-element group 22: 	 branch_block_stmt_31/assign_stmt_52_to_assign_stmt_70/slice_65_update_start_
      -- CP-element group 22: 	 branch_block_stmt_31/assign_stmt_52_to_assign_stmt_70/slice_65_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_31/assign_stmt_52_to_assign_stmt_70/R_head1_63_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_31/assign_stmt_52_to_assign_stmt_70/R_head1_63_sample_completed_
      -- CP-element group 22: 	 branch_block_stmt_31/assign_stmt_52_to_assign_stmt_70/R_head1_63_update_start_
      -- CP-element group 22: 	 branch_block_stmt_31/assign_stmt_52_to_assign_stmt_70/R_head1_63_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_31/assign_stmt_52_to_assign_stmt_70/slice_65_Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_31/assign_stmt_52_to_assign_stmt_70/slice_65_Sample/$exit
      -- CP-element group 22: 	 branch_block_stmt_31/assign_stmt_52_to_assign_stmt_70/slice_65_Sample/rr
      -- CP-element group 22: 	 branch_block_stmt_31/assign_stmt_52_to_assign_stmt_70/slice_65_Sample/ra
      -- CP-element group 22: 	 branch_block_stmt_31/assign_stmt_52_to_assign_stmt_70/slice_65_Update/$entry
      -- CP-element group 22: 	 branch_block_stmt_31/assign_stmt_52_to_assign_stmt_70/slice_65_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_31/assign_stmt_52_to_assign_stmt_70/slice_65_Update/cr
      -- CP-element group 22: 	 branch_block_stmt_31/assign_stmt_52_to_assign_stmt_70/slice_65_Update/ca
      -- CP-element group 22: 	 branch_block_stmt_31/assign_stmt_52_to_assign_stmt_70/slice_69_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_31/assign_stmt_52_to_assign_stmt_70/slice_69_sample_completed_
      -- CP-element group 22: 	 branch_block_stmt_31/assign_stmt_52_to_assign_stmt_70/slice_69_update_start_
      -- CP-element group 22: 	 branch_block_stmt_31/assign_stmt_52_to_assign_stmt_70/slice_69_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_31/assign_stmt_52_to_assign_stmt_70/R_head1_68_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_31/assign_stmt_52_to_assign_stmt_70/R_head1_68_sample_completed_
      -- CP-element group 22: 	 branch_block_stmt_31/assign_stmt_52_to_assign_stmt_70/R_head1_68_update_start_
      -- CP-element group 22: 	 branch_block_stmt_31/assign_stmt_52_to_assign_stmt_70/R_head1_68_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_31/assign_stmt_52_to_assign_stmt_70/slice_69_Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_31/assign_stmt_52_to_assign_stmt_70/slice_69_Sample/$exit
      -- CP-element group 22: 	 branch_block_stmt_31/assign_stmt_52_to_assign_stmt_70/slice_69_Sample/rr
      -- CP-element group 22: 	 branch_block_stmt_31/assign_stmt_52_to_assign_stmt_70/slice_69_Sample/ra
      -- CP-element group 22: 	 branch_block_stmt_31/assign_stmt_52_to_assign_stmt_70/slice_69_Update/$entry
      -- CP-element group 22: 	 branch_block_stmt_31/assign_stmt_52_to_assign_stmt_70/slice_69_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_31/assign_stmt_52_to_assign_stmt_70/slice_69_Update/cr
      -- CP-element group 22: 	 branch_block_stmt_31/assign_stmt_52_to_assign_stmt_70/slice_69_Update/ca
      -- 
    In_wrap_daemon_CP_0_elements(22) <= In_wrap_daemon_CP_0_elements(5);
    -- CP-element group 23:  transition  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	6 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (1) 
      -- CP-element group 23: 	 branch_block_stmt_31/if_stmt_71_dead_link/$entry
      -- 
    In_wrap_daemon_CP_0_elements(23) <= In_wrap_daemon_CP_0_elements(6);
    -- CP-element group 24:  transition  output  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	6 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24:  members (17) 
      -- CP-element group 24: 	 branch_block_stmt_31/if_stmt_71_eval_test/$entry
      -- CP-element group 24: 	 branch_block_stmt_31/if_stmt_71_eval_test/$exit
      -- CP-element group 24: 	 branch_block_stmt_31/if_stmt_71_eval_test/EQ_u1_u1_74/$entry
      -- CP-element group 24: 	 branch_block_stmt_31/if_stmt_71_eval_test/EQ_u1_u1_74/$exit
      -- CP-element group 24: 	 branch_block_stmt_31/if_stmt_71_eval_test/EQ_u1_u1_74/EQ_u1_u1_74_inputs/$entry
      -- CP-element group 24: 	 branch_block_stmt_31/if_stmt_71_eval_test/EQ_u1_u1_74/EQ_u1_u1_74_inputs/$exit
      -- CP-element group 24: 	 branch_block_stmt_31/if_stmt_71_eval_test/EQ_u1_u1_74/SplitProtocol/$entry
      -- CP-element group 24: 	 branch_block_stmt_31/if_stmt_71_eval_test/EQ_u1_u1_74/SplitProtocol/$exit
      -- CP-element group 24: 	 branch_block_stmt_31/if_stmt_71_eval_test/EQ_u1_u1_74/SplitProtocol/Sample/$entry
      -- CP-element group 24: 	 branch_block_stmt_31/if_stmt_71_eval_test/EQ_u1_u1_74/SplitProtocol/Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_31/if_stmt_71_eval_test/EQ_u1_u1_74/SplitProtocol/Sample/rr
      -- CP-element group 24: 	 branch_block_stmt_31/if_stmt_71_eval_test/EQ_u1_u1_74/SplitProtocol/Sample/ra
      -- CP-element group 24: 	 branch_block_stmt_31/if_stmt_71_eval_test/EQ_u1_u1_74/SplitProtocol/Update/$entry
      -- CP-element group 24: 	 branch_block_stmt_31/if_stmt_71_eval_test/EQ_u1_u1_74/SplitProtocol/Update/$exit
      -- CP-element group 24: 	 branch_block_stmt_31/if_stmt_71_eval_test/EQ_u1_u1_74/SplitProtocol/Update/cr
      -- CP-element group 24: 	 branch_block_stmt_31/if_stmt_71_eval_test/EQ_u1_u1_74/SplitProtocol/Update/ca
      -- CP-element group 24: 	 branch_block_stmt_31/if_stmt_71_eval_test/branch_req
      -- 
    branch_req_247_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_247_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => In_wrap_daemon_CP_0_elements(24), ack => if_stmt_71_branch_req_0); -- 
    In_wrap_daemon_CP_0_elements(24) <= In_wrap_daemon_CP_0_elements(6);
    -- CP-element group 25:  branch  place  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	24 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25: 	28 
    -- CP-element group 25:  members (1) 
      -- CP-element group 25: 	 branch_block_stmt_31/EQ_u1_u1_74_place
      -- 
    In_wrap_daemon_CP_0_elements(25) <= In_wrap_daemon_CP_0_elements(24);
    -- CP-element group 26:  transition  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	25 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	27 
    -- CP-element group 26:  members (1) 
      -- CP-element group 26: 	 branch_block_stmt_31/if_stmt_71_if_link/$entry
      -- 
    In_wrap_daemon_CP_0_elements(26) <= In_wrap_daemon_CP_0_elements(25);
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	26 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	30 
    -- CP-element group 27:  members (2) 
      -- CP-element group 27: 	 branch_block_stmt_31/if_stmt_71_if_link/$exit
      -- CP-element group 27: 	 branch_block_stmt_31/if_stmt_71_if_link/if_choice_transition
      -- 
    if_choice_transition_252_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_71_branch_ack_1, ack => In_wrap_daemon_CP_0_elements(27)); -- 
    -- CP-element group 28:  transition  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	25 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28:  members (1) 
      -- CP-element group 28: 	 branch_block_stmt_31/if_stmt_71_else_link/$entry
      -- 
    In_wrap_daemon_CP_0_elements(28) <= In_wrap_daemon_CP_0_elements(25);
    -- CP-element group 29:  transition  input  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	28 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	7 
    -- CP-element group 29:  members (2) 
      -- CP-element group 29: 	 branch_block_stmt_31/if_stmt_71_else_link/$exit
      -- CP-element group 29: 	 branch_block_stmt_31/if_stmt_71_else_link/else_choice_transition
      -- 
    else_choice_transition_256_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_71_branch_ack_0, ack => In_wrap_daemon_CP_0_elements(29)); -- 
    -- CP-element group 30:  place  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	27 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	35 
    -- CP-element group 30:  members (1) 
      -- CP-element group 30: 	 branch_block_stmt_31/assign_stmt_77__entry__
      -- 
    In_wrap_daemon_CP_0_elements(30) <= In_wrap_daemon_CP_0_elements(27);
    -- CP-element group 31:  place  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	37 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	38 
    -- CP-element group 31:  members (2) 
      -- CP-element group 31: 	 branch_block_stmt_31/assign_stmt_77__exit__
      -- CP-element group 31: 	 branch_block_stmt_31/assign_stmt_81_to_assign_stmt_85__entry__
      -- 
    In_wrap_daemon_CP_0_elements(31) <= In_wrap_daemon_CP_0_elements(37);
    -- CP-element group 32:  place  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	43 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	44 
    -- CP-element group 32:  members (2) 
      -- CP-element group 32: 	 branch_block_stmt_31/assign_stmt_81_to_assign_stmt_85__exit__
      -- CP-element group 32: 	 branch_block_stmt_31/assign_stmt_88__entry__
      -- 
    In_wrap_daemon_CP_0_elements(32) <= In_wrap_daemon_CP_0_elements(43);
    -- CP-element group 33:  place  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	46 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	47 
    -- CP-element group 33:  members (2) 
      -- CP-element group 33: 	 branch_block_stmt_31/assign_stmt_88__exit__
      -- CP-element group 33: 	 branch_block_stmt_31/assign_stmt_91__entry__
      -- 
    In_wrap_daemon_CP_0_elements(33) <= In_wrap_daemon_CP_0_elements(46);
    -- CP-element group 34:  place  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	49 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	7 
    -- CP-element group 34:  members (1) 
      -- CP-element group 34: 	 branch_block_stmt_31/assign_stmt_91__exit__
      -- 
    In_wrap_daemon_CP_0_elements(34) <= In_wrap_daemon_CP_0_elements(49);
    -- CP-element group 35:  transition  output  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	30 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	36 
    -- CP-element group 35:  members (4) 
      -- CP-element group 35: 	 branch_block_stmt_31/assign_stmt_77/$entry
      -- CP-element group 35: 	 branch_block_stmt_31/assign_stmt_77/RPIPE_w_in_buf_76_sample_start_
      -- CP-element group 35: 	 branch_block_stmt_31/assign_stmt_77/RPIPE_w_in_buf_76_Sample/$entry
      -- CP-element group 35: 	 branch_block_stmt_31/assign_stmt_77/RPIPE_w_in_buf_76_Sample/rr
      -- 
    rr_275_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_275_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => In_wrap_daemon_CP_0_elements(35), ack => RPIPE_w_in_buf_76_inst_req_0); -- 
    In_wrap_daemon_CP_0_elements(35) <= In_wrap_daemon_CP_0_elements(30);
    -- CP-element group 36:  transition  input  output  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	35 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	37 
    -- CP-element group 36:  members (6) 
      -- CP-element group 36: 	 branch_block_stmt_31/assign_stmt_77/RPIPE_w_in_buf_76_sample_completed_
      -- CP-element group 36: 	 branch_block_stmt_31/assign_stmt_77/RPIPE_w_in_buf_76_update_start_
      -- CP-element group 36: 	 branch_block_stmt_31/assign_stmt_77/RPIPE_w_in_buf_76_Sample/$exit
      -- CP-element group 36: 	 branch_block_stmt_31/assign_stmt_77/RPIPE_w_in_buf_76_Sample/ra
      -- CP-element group 36: 	 branch_block_stmt_31/assign_stmt_77/RPIPE_w_in_buf_76_Update/$entry
      -- CP-element group 36: 	 branch_block_stmt_31/assign_stmt_77/RPIPE_w_in_buf_76_Update/cr
      -- 
    ra_276_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_w_in_buf_76_inst_ack_0, ack => In_wrap_daemon_CP_0_elements(36)); -- 
    cr_280_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_280_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => In_wrap_daemon_CP_0_elements(36), ack => RPIPE_w_in_buf_76_inst_req_1); -- 
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	36 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	31 
    -- CP-element group 37:  members (4) 
      -- CP-element group 37: 	 branch_block_stmt_31/assign_stmt_77/$exit
      -- CP-element group 37: 	 branch_block_stmt_31/assign_stmt_77/RPIPE_w_in_buf_76_update_completed_
      -- CP-element group 37: 	 branch_block_stmt_31/assign_stmt_77/RPIPE_w_in_buf_76_Update/$exit
      -- CP-element group 37: 	 branch_block_stmt_31/assign_stmt_77/RPIPE_w_in_buf_76_Update/ca
      -- 
    ca_281_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_w_in_buf_76_inst_ack_1, ack => In_wrap_daemon_CP_0_elements(37)); -- 
    -- CP-element group 38:  fork  transition  output  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	31 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38: 	40 
    -- CP-element group 38: 	41 
    -- CP-element group 38: 	42 
    -- CP-element group 38:  members (21) 
      -- CP-element group 38: 	 branch_block_stmt_31/assign_stmt_81_to_assign_stmt_85/$entry
      -- CP-element group 38: 	 branch_block_stmt_31/assign_stmt_81_to_assign_stmt_85/slice_80_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_31/assign_stmt_81_to_assign_stmt_85/slice_80_update_start_
      -- CP-element group 38: 	 branch_block_stmt_31/assign_stmt_81_to_assign_stmt_85/R_key_79_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_31/assign_stmt_81_to_assign_stmt_85/R_key_79_sample_completed_
      -- CP-element group 38: 	 branch_block_stmt_31/assign_stmt_81_to_assign_stmt_85/R_key_79_update_start_
      -- CP-element group 38: 	 branch_block_stmt_31/assign_stmt_81_to_assign_stmt_85/R_key_79_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_31/assign_stmt_81_to_assign_stmt_85/slice_80_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_31/assign_stmt_81_to_assign_stmt_85/slice_80_Sample/rr
      -- CP-element group 38: 	 branch_block_stmt_31/assign_stmt_81_to_assign_stmt_85/slice_80_Update/$entry
      -- CP-element group 38: 	 branch_block_stmt_31/assign_stmt_81_to_assign_stmt_85/slice_80_Update/cr
      -- CP-element group 38: 	 branch_block_stmt_31/assign_stmt_81_to_assign_stmt_85/slice_84_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_31/assign_stmt_81_to_assign_stmt_85/slice_84_update_start_
      -- CP-element group 38: 	 branch_block_stmt_31/assign_stmt_81_to_assign_stmt_85/R_key_83_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_31/assign_stmt_81_to_assign_stmt_85/R_key_83_sample_completed_
      -- CP-element group 38: 	 branch_block_stmt_31/assign_stmt_81_to_assign_stmt_85/R_key_83_update_start_
      -- CP-element group 38: 	 branch_block_stmt_31/assign_stmt_81_to_assign_stmt_85/R_key_83_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_31/assign_stmt_81_to_assign_stmt_85/slice_84_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_31/assign_stmt_81_to_assign_stmt_85/slice_84_Sample/rr
      -- CP-element group 38: 	 branch_block_stmt_31/assign_stmt_81_to_assign_stmt_85/slice_84_Update/$entry
      -- CP-element group 38: 	 branch_block_stmt_31/assign_stmt_81_to_assign_stmt_85/slice_84_Update/cr
      -- 
    cr_301_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_301_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => In_wrap_daemon_CP_0_elements(38), ack => slice_80_inst_req_1); -- 
    rr_296_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_296_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => In_wrap_daemon_CP_0_elements(38), ack => slice_80_inst_req_0); -- 
    cr_319_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_319_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => In_wrap_daemon_CP_0_elements(38), ack => slice_84_inst_req_1); -- 
    rr_314_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_314_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => In_wrap_daemon_CP_0_elements(38), ack => slice_84_inst_req_0); -- 
    In_wrap_daemon_CP_0_elements(38) <= In_wrap_daemon_CP_0_elements(31);
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_31/assign_stmt_81_to_assign_stmt_85/slice_80_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_31/assign_stmt_81_to_assign_stmt_85/slice_80_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_31/assign_stmt_81_to_assign_stmt_85/slice_80_Sample/ra
      -- 
    ra_297_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_80_inst_ack_0, ack => In_wrap_daemon_CP_0_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	38 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	43 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_31/assign_stmt_81_to_assign_stmt_85/slice_80_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_31/assign_stmt_81_to_assign_stmt_85/slice_80_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_31/assign_stmt_81_to_assign_stmt_85/slice_80_Update/ca
      -- 
    ca_302_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_80_inst_ack_1, ack => In_wrap_daemon_CP_0_elements(40)); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	38 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_31/assign_stmt_81_to_assign_stmt_85/slice_84_sample_completed_
      -- CP-element group 41: 	 branch_block_stmt_31/assign_stmt_81_to_assign_stmt_85/slice_84_Sample/$exit
      -- CP-element group 41: 	 branch_block_stmt_31/assign_stmt_81_to_assign_stmt_85/slice_84_Sample/ra
      -- 
    ra_315_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_84_inst_ack_0, ack => In_wrap_daemon_CP_0_elements(41)); -- 
    -- CP-element group 42:  transition  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	38 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_31/assign_stmt_81_to_assign_stmt_85/slice_84_update_completed_
      -- CP-element group 42: 	 branch_block_stmt_31/assign_stmt_81_to_assign_stmt_85/slice_84_Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_31/assign_stmt_81_to_assign_stmt_85/slice_84_Update/ca
      -- 
    ca_320_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_84_inst_ack_1, ack => In_wrap_daemon_CP_0_elements(42)); -- 
    -- CP-element group 43:  join  transition  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	40 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	32 
    -- CP-element group 43:  members (1) 
      -- CP-element group 43: 	 branch_block_stmt_31/assign_stmt_81_to_assign_stmt_85/$exit
      -- 
    In_wrap_daemon_cp_element_group_43: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "In_wrap_daemon_cp_element_group_43"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= In_wrap_daemon_CP_0_elements(40) & In_wrap_daemon_CP_0_elements(42);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => In_wrap_daemon_CP_0_elements(43), clk => clk, reset => reset); --
    end block;
    -- CP-element group 44:  transition  output  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	32 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	45 
    -- CP-element group 44:  members (8) 
      -- CP-element group 44: 	 branch_block_stmt_31/assign_stmt_88/$entry
      -- CP-element group 44: 	 branch_block_stmt_31/assign_stmt_88/R_keyA_87_sample_start_
      -- CP-element group 44: 	 branch_block_stmt_31/assign_stmt_88/R_keyA_87_sample_completed_
      -- CP-element group 44: 	 branch_block_stmt_31/assign_stmt_88/R_keyA_87_update_start_
      -- CP-element group 44: 	 branch_block_stmt_31/assign_stmt_88/R_keyA_87_update_completed_
      -- CP-element group 44: 	 branch_block_stmt_31/assign_stmt_88/WPIPE_cmd_in_86_sample_start_
      -- CP-element group 44: 	 branch_block_stmt_31/assign_stmt_88/WPIPE_cmd_in_86_Sample/$entry
      -- CP-element group 44: 	 branch_block_stmt_31/assign_stmt_88/WPIPE_cmd_in_86_Sample/req
      -- 
    req_335_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_335_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => In_wrap_daemon_CP_0_elements(44), ack => WPIPE_cmd_in_86_inst_req_0); -- 
    In_wrap_daemon_CP_0_elements(44) <= In_wrap_daemon_CP_0_elements(32);
    -- CP-element group 45:  transition  input  output  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	44 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45:  members (6) 
      -- CP-element group 45: 	 branch_block_stmt_31/assign_stmt_88/WPIPE_cmd_in_86_sample_completed_
      -- CP-element group 45: 	 branch_block_stmt_31/assign_stmt_88/WPIPE_cmd_in_86_update_start_
      -- CP-element group 45: 	 branch_block_stmt_31/assign_stmt_88/WPIPE_cmd_in_86_Sample/$exit
      -- CP-element group 45: 	 branch_block_stmt_31/assign_stmt_88/WPIPE_cmd_in_86_Sample/ack
      -- CP-element group 45: 	 branch_block_stmt_31/assign_stmt_88/WPIPE_cmd_in_86_Update/$entry
      -- CP-element group 45: 	 branch_block_stmt_31/assign_stmt_88/WPIPE_cmd_in_86_Update/req
      -- 
    ack_336_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_cmd_in_86_inst_ack_0, ack => In_wrap_daemon_CP_0_elements(45)); -- 
    req_340_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_340_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => In_wrap_daemon_CP_0_elements(45), ack => WPIPE_cmd_in_86_inst_req_1); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	33 
    -- CP-element group 46:  members (4) 
      -- CP-element group 46: 	 branch_block_stmt_31/assign_stmt_88/$exit
      -- CP-element group 46: 	 branch_block_stmt_31/assign_stmt_88/WPIPE_cmd_in_86_update_completed_
      -- CP-element group 46: 	 branch_block_stmt_31/assign_stmt_88/WPIPE_cmd_in_86_Update/$exit
      -- CP-element group 46: 	 branch_block_stmt_31/assign_stmt_88/WPIPE_cmd_in_86_Update/ack
      -- 
    ack_341_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_cmd_in_86_inst_ack_1, ack => In_wrap_daemon_CP_0_elements(46)); -- 
    -- CP-element group 47:  transition  output  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	33 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	48 
    -- CP-element group 47:  members (8) 
      -- CP-element group 47: 	 branch_block_stmt_31/assign_stmt_91/WPIPE_cmd_in_89_Sample/$entry
      -- CP-element group 47: 	 branch_block_stmt_31/assign_stmt_91/WPIPE_cmd_in_89_Sample/req
      -- CP-element group 47: 	 branch_block_stmt_31/assign_stmt_91/$entry
      -- CP-element group 47: 	 branch_block_stmt_31/assign_stmt_91/R_keyB_90_sample_start_
      -- CP-element group 47: 	 branch_block_stmt_31/assign_stmt_91/R_keyB_90_sample_completed_
      -- CP-element group 47: 	 branch_block_stmt_31/assign_stmt_91/R_keyB_90_update_start_
      -- CP-element group 47: 	 branch_block_stmt_31/assign_stmt_91/R_keyB_90_update_completed_
      -- CP-element group 47: 	 branch_block_stmt_31/assign_stmt_91/WPIPE_cmd_in_89_sample_start_
      -- 
    req_356_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_356_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => In_wrap_daemon_CP_0_elements(47), ack => WPIPE_cmd_in_89_inst_req_0); -- 
    In_wrap_daemon_CP_0_elements(47) <= In_wrap_daemon_CP_0_elements(33);
    -- CP-element group 48:  transition  input  output  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	47 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	49 
    -- CP-element group 48:  members (6) 
      -- CP-element group 48: 	 branch_block_stmt_31/assign_stmt_91/WPIPE_cmd_in_89_sample_completed_
      -- CP-element group 48: 	 branch_block_stmt_31/assign_stmt_91/WPIPE_cmd_in_89_update_start_
      -- CP-element group 48: 	 branch_block_stmt_31/assign_stmt_91/WPIPE_cmd_in_89_Sample/$exit
      -- CP-element group 48: 	 branch_block_stmt_31/assign_stmt_91/WPIPE_cmd_in_89_Sample/ack
      -- CP-element group 48: 	 branch_block_stmt_31/assign_stmt_91/WPIPE_cmd_in_89_Update/$entry
      -- CP-element group 48: 	 branch_block_stmt_31/assign_stmt_91/WPIPE_cmd_in_89_Update/req
      -- 
    ack_357_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_cmd_in_89_inst_ack_0, ack => In_wrap_daemon_CP_0_elements(48)); -- 
    req_361_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_361_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => In_wrap_daemon_CP_0_elements(48), ack => WPIPE_cmd_in_89_inst_req_1); -- 
    -- CP-element group 49:  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	48 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	34 
    -- CP-element group 49:  members (4) 
      -- CP-element group 49: 	 branch_block_stmt_31/assign_stmt_91/WPIPE_cmd_in_89_update_completed_
      -- CP-element group 49: 	 branch_block_stmt_31/assign_stmt_91/WPIPE_cmd_in_89_Update/$exit
      -- CP-element group 49: 	 branch_block_stmt_31/assign_stmt_91/WPIPE_cmd_in_89_Update/ack
      -- CP-element group 49: 	 branch_block_stmt_31/assign_stmt_91/$exit
      -- 
    ack_362_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_cmd_in_89_inst_ack_1, ack => In_wrap_daemon_CP_0_elements(49)); -- 
    -- CP-element group 50:  join  fork  transition  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	7 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50: 	52 
    -- CP-element group 50:  members (67) 
      -- CP-element group 50: 	 branch_block_stmt_31/assign_stmt_107/$entry
      -- CP-element group 50: 	 branch_block_stmt_31/assign_stmt_107/OR_u15_u15_106_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_31/assign_stmt_107/OR_u15_u15_106_update_start_
      -- CP-element group 50: 	 branch_block_stmt_31/assign_stmt_107/MUX_99_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_31/assign_stmt_107/MUX_99_sample_completed_
      -- CP-element group 50: 	 branch_block_stmt_31/assign_stmt_107/MUX_99_update_start_
      -- CP-element group 50: 	 branch_block_stmt_31/assign_stmt_107/MUX_99_update_completed_
      -- CP-element group 50: 	 branch_block_stmt_31/assign_stmt_107/ULT_u15_u1_96_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_31/assign_stmt_107/ULT_u15_u1_96_sample_completed_
      -- CP-element group 50: 	 branch_block_stmt_31/assign_stmt_107/ULT_u15_u1_96_update_start_
      -- CP-element group 50: 	 branch_block_stmt_31/assign_stmt_107/ULT_u15_u1_96_update_completed_
      -- CP-element group 50: 	 branch_block_stmt_31/assign_stmt_107/R_count_95_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_31/assign_stmt_107/R_count_95_sample_completed_
      -- CP-element group 50: 	 branch_block_stmt_31/assign_stmt_107/R_count_95_update_start_
      -- CP-element group 50: 	 branch_block_stmt_31/assign_stmt_107/R_count_95_update_completed_
      -- CP-element group 50: 	 branch_block_stmt_31/assign_stmt_107/ULT_u15_u1_96_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_31/assign_stmt_107/ULT_u15_u1_96_Sample/$exit
      -- CP-element group 50: 	 branch_block_stmt_31/assign_stmt_107/ULT_u15_u1_96_Sample/rr
      -- CP-element group 50: 	 branch_block_stmt_31/assign_stmt_107/ULT_u15_u1_96_Sample/ra
      -- CP-element group 50: 	 branch_block_stmt_31/assign_stmt_107/ULT_u15_u1_96_Update/$entry
      -- CP-element group 50: 	 branch_block_stmt_31/assign_stmt_107/ULT_u15_u1_96_Update/$exit
      -- CP-element group 50: 	 branch_block_stmt_31/assign_stmt_107/ULT_u15_u1_96_Update/cr
      -- CP-element group 50: 	 branch_block_stmt_31/assign_stmt_107/ULT_u15_u1_96_Update/ca
      -- CP-element group 50: 	 branch_block_stmt_31/assign_stmt_107/MUX_99_start/$entry
      -- CP-element group 50: 	 branch_block_stmt_31/assign_stmt_107/MUX_99_start/$exit
      -- CP-element group 50: 	 branch_block_stmt_31/assign_stmt_107/MUX_99_start/req
      -- CP-element group 50: 	 branch_block_stmt_31/assign_stmt_107/MUX_99_start/ack
      -- CP-element group 50: 	 branch_block_stmt_31/assign_stmt_107/MUX_99_complete/$entry
      -- CP-element group 50: 	 branch_block_stmt_31/assign_stmt_107/MUX_99_complete/$exit
      -- CP-element group 50: 	 branch_block_stmt_31/assign_stmt_107/MUX_99_complete/req
      -- CP-element group 50: 	 branch_block_stmt_31/assign_stmt_107/MUX_99_complete/ack
      -- CP-element group 50: 	 branch_block_stmt_31/assign_stmt_107/MUX_105_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_31/assign_stmt_107/MUX_105_sample_completed_
      -- CP-element group 50: 	 branch_block_stmt_31/assign_stmt_107/MUX_105_update_start_
      -- CP-element group 50: 	 branch_block_stmt_31/assign_stmt_107/MUX_105_update_completed_
      -- CP-element group 50: 	 branch_block_stmt_31/assign_stmt_107/UGE_u15_u1_102_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_31/assign_stmt_107/UGE_u15_u1_102_sample_completed_
      -- CP-element group 50: 	 branch_block_stmt_31/assign_stmt_107/UGE_u15_u1_102_update_start_
      -- CP-element group 50: 	 branch_block_stmt_31/assign_stmt_107/UGE_u15_u1_102_update_completed_
      -- CP-element group 50: 	 branch_block_stmt_31/assign_stmt_107/R_count_101_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_31/assign_stmt_107/R_count_101_sample_completed_
      -- CP-element group 50: 	 branch_block_stmt_31/assign_stmt_107/R_count_101_update_start_
      -- CP-element group 50: 	 branch_block_stmt_31/assign_stmt_107/R_count_101_update_completed_
      -- CP-element group 50: 	 branch_block_stmt_31/assign_stmt_107/UGE_u15_u1_102_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_31/assign_stmt_107/UGE_u15_u1_102_Sample/$exit
      -- CP-element group 50: 	 branch_block_stmt_31/assign_stmt_107/UGE_u15_u1_102_Sample/rr
      -- CP-element group 50: 	 branch_block_stmt_31/assign_stmt_107/UGE_u15_u1_102_Sample/ra
      -- CP-element group 50: 	 branch_block_stmt_31/assign_stmt_107/UGE_u15_u1_102_Update/$entry
      -- CP-element group 50: 	 branch_block_stmt_31/assign_stmt_107/UGE_u15_u1_102_Update/$exit
      -- CP-element group 50: 	 branch_block_stmt_31/assign_stmt_107/UGE_u15_u1_102_Update/cr
      -- CP-element group 50: 	 branch_block_stmt_31/assign_stmt_107/UGE_u15_u1_102_Update/ca
      -- CP-element group 50: 	 branch_block_stmt_31/assign_stmt_107/R_count_103_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_31/assign_stmt_107/R_count_103_sample_completed_
      -- CP-element group 50: 	 branch_block_stmt_31/assign_stmt_107/R_count_103_update_start_
      -- CP-element group 50: 	 branch_block_stmt_31/assign_stmt_107/R_count_103_update_completed_
      -- CP-element group 50: 	 branch_block_stmt_31/assign_stmt_107/MUX_105_start/$entry
      -- CP-element group 50: 	 branch_block_stmt_31/assign_stmt_107/MUX_105_start/$exit
      -- CP-element group 50: 	 branch_block_stmt_31/assign_stmt_107/MUX_105_start/req
      -- CP-element group 50: 	 branch_block_stmt_31/assign_stmt_107/MUX_105_start/ack
      -- CP-element group 50: 	 branch_block_stmt_31/assign_stmt_107/MUX_105_complete/$entry
      -- CP-element group 50: 	 branch_block_stmt_31/assign_stmt_107/MUX_105_complete/$exit
      -- CP-element group 50: 	 branch_block_stmt_31/assign_stmt_107/MUX_105_complete/req
      -- CP-element group 50: 	 branch_block_stmt_31/assign_stmt_107/MUX_105_complete/ack
      -- CP-element group 50: 	 branch_block_stmt_31/assign_stmt_107/OR_u15_u15_106_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_31/assign_stmt_107/OR_u15_u15_106_Sample/rr
      -- CP-element group 50: 	 branch_block_stmt_31/assign_stmt_107/OR_u15_u15_106_Update/$entry
      -- CP-element group 50: 	 branch_block_stmt_31/assign_stmt_107/OR_u15_u15_106_Update/cr
      -- 
    cr_446_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_446_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => In_wrap_daemon_CP_0_elements(50), ack => OR_u15_u15_106_inst_req_1); -- 
    rr_441_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_441_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => In_wrap_daemon_CP_0_elements(50), ack => OR_u15_u15_106_inst_req_0); -- 
    In_wrap_daemon_CP_0_elements(50) <= In_wrap_daemon_CP_0_elements(7);
    -- CP-element group 51:  transition  input  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 branch_block_stmt_31/assign_stmt_107/OR_u15_u15_106_sample_completed_
      -- CP-element group 51: 	 branch_block_stmt_31/assign_stmt_107/OR_u15_u15_106_Sample/$exit
      -- CP-element group 51: 	 branch_block_stmt_31/assign_stmt_107/OR_u15_u15_106_Sample/ra
      -- 
    ra_442_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => OR_u15_u15_106_inst_ack_0, ack => In_wrap_daemon_CP_0_elements(51)); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	50 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	8 
    -- CP-element group 52:  members (4) 
      -- CP-element group 52: 	 branch_block_stmt_31/assign_stmt_107/$exit
      -- CP-element group 52: 	 branch_block_stmt_31/assign_stmt_107/OR_u15_u15_106_update_completed_
      -- CP-element group 52: 	 branch_block_stmt_31/assign_stmt_107/OR_u15_u15_106_Update/$exit
      -- CP-element group 52: 	 branch_block_stmt_31/assign_stmt_107/OR_u15_u15_106_Update/ca
      -- 
    ca_447_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => OR_u15_u15_106_inst_ack_1, ack => In_wrap_daemon_CP_0_elements(52)); -- 
    -- CP-element group 53:  transition  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	9 
    -- CP-element group 53: successors 
    -- CP-element group 53:  members (1) 
      -- CP-element group 53: 	 branch_block_stmt_31/if_stmt_114_dead_link/$entry
      -- 
    In_wrap_daemon_CP_0_elements(53) <= In_wrap_daemon_CP_0_elements(9);
    -- CP-element group 54:  transition  output  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	9 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	55 
    -- CP-element group 54:  members (17) 
      -- CP-element group 54: 	 branch_block_stmt_31/if_stmt_114_eval_test/$entry
      -- CP-element group 54: 	 branch_block_stmt_31/if_stmt_114_eval_test/$exit
      -- CP-element group 54: 	 branch_block_stmt_31/if_stmt_114_eval_test/EQ_u1_u1_117/$entry
      -- CP-element group 54: 	 branch_block_stmt_31/if_stmt_114_eval_test/EQ_u1_u1_117/$exit
      -- CP-element group 54: 	 branch_block_stmt_31/if_stmt_114_eval_test/EQ_u1_u1_117/EQ_u1_u1_117_inputs/$entry
      -- CP-element group 54: 	 branch_block_stmt_31/if_stmt_114_eval_test/EQ_u1_u1_117/EQ_u1_u1_117_inputs/$exit
      -- CP-element group 54: 	 branch_block_stmt_31/if_stmt_114_eval_test/EQ_u1_u1_117/SplitProtocol/$entry
      -- CP-element group 54: 	 branch_block_stmt_31/if_stmt_114_eval_test/EQ_u1_u1_117/SplitProtocol/$exit
      -- CP-element group 54: 	 branch_block_stmt_31/if_stmt_114_eval_test/EQ_u1_u1_117/SplitProtocol/Sample/$entry
      -- CP-element group 54: 	 branch_block_stmt_31/if_stmt_114_eval_test/EQ_u1_u1_117/SplitProtocol/Sample/$exit
      -- CP-element group 54: 	 branch_block_stmt_31/if_stmt_114_eval_test/EQ_u1_u1_117/SplitProtocol/Sample/rr
      -- CP-element group 54: 	 branch_block_stmt_31/if_stmt_114_eval_test/EQ_u1_u1_117/SplitProtocol/Sample/ra
      -- CP-element group 54: 	 branch_block_stmt_31/if_stmt_114_eval_test/EQ_u1_u1_117/SplitProtocol/Update/$entry
      -- CP-element group 54: 	 branch_block_stmt_31/if_stmt_114_eval_test/EQ_u1_u1_117/SplitProtocol/Update/$exit
      -- CP-element group 54: 	 branch_block_stmt_31/if_stmt_114_eval_test/EQ_u1_u1_117/SplitProtocol/Update/cr
      -- CP-element group 54: 	 branch_block_stmt_31/if_stmt_114_eval_test/EQ_u1_u1_117/SplitProtocol/Update/ca
      -- CP-element group 54: 	 branch_block_stmt_31/if_stmt_114_eval_test/branch_req
      -- 
    branch_req_474_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_474_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => In_wrap_daemon_CP_0_elements(54), ack => if_stmt_114_branch_req_0); -- 
    In_wrap_daemon_CP_0_elements(54) <= In_wrap_daemon_CP_0_elements(9);
    -- CP-element group 55:  branch  place  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	54 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55: 	58 
    -- CP-element group 55:  members (1) 
      -- CP-element group 55: 	 branch_block_stmt_31/EQ_u1_u1_117_place
      -- 
    In_wrap_daemon_CP_0_elements(55) <= In_wrap_daemon_CP_0_elements(54);
    -- CP-element group 56:  transition  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	57 
    -- CP-element group 56:  members (1) 
      -- CP-element group 56: 	 branch_block_stmt_31/if_stmt_114_if_link/$entry
      -- 
    In_wrap_daemon_CP_0_elements(56) <= In_wrap_daemon_CP_0_elements(55);
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	56 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	60 
    -- CP-element group 57:  members (2) 
      -- CP-element group 57: 	 branch_block_stmt_31/if_stmt_114_if_link/$exit
      -- CP-element group 57: 	 branch_block_stmt_31/if_stmt_114_if_link/if_choice_transition
      -- 
    if_choice_transition_479_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_114_branch_ack_1, ack => In_wrap_daemon_CP_0_elements(57)); -- 
    -- CP-element group 58:  transition  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	55 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58:  members (1) 
      -- CP-element group 58: 	 branch_block_stmt_31/if_stmt_114_else_link/$entry
      -- 
    In_wrap_daemon_CP_0_elements(58) <= In_wrap_daemon_CP_0_elements(55);
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	67 
    -- CP-element group 59:  members (2) 
      -- CP-element group 59: 	 branch_block_stmt_31/if_stmt_114_else_link/$exit
      -- CP-element group 59: 	 branch_block_stmt_31/if_stmt_114_else_link/else_choice_transition
      -- 
    else_choice_transition_483_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_114_branch_ack_0, ack => In_wrap_daemon_CP_0_elements(59)); -- 
    -- CP-element group 60:  place  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	57 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	62 
    -- CP-element group 60:  members (1) 
      -- CP-element group 60: 	 branch_block_stmt_31/assign_stmt_120__entry__
      -- 
    In_wrap_daemon_CP_0_elements(60) <= In_wrap_daemon_CP_0_elements(57);
    -- CP-element group 61:  place  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	66 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	10 
    -- CP-element group 61:  members (1) 
      -- CP-element group 61: 	 branch_block_stmt_31/assign_stmt_120__exit__
      -- 
    In_wrap_daemon_CP_0_elements(61) <= In_wrap_daemon_CP_0_elements(66);
    -- CP-element group 62:  transition  output  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	60 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62:  members (4) 
      -- CP-element group 62: 	 branch_block_stmt_31/assign_stmt_120/$entry
      -- CP-element group 62: 	 branch_block_stmt_31/assign_stmt_120/RPIPE_w_in_buf_119_sample_start_
      -- CP-element group 62: 	 branch_block_stmt_31/assign_stmt_120/RPIPE_w_in_buf_119_Sample/$entry
      -- CP-element group 62: 	 branch_block_stmt_31/assign_stmt_120/RPIPE_w_in_buf_119_Sample/rr
      -- 
    rr_496_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_496_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => In_wrap_daemon_CP_0_elements(62), ack => RPIPE_w_in_buf_119_inst_req_0); -- 
    In_wrap_daemon_CP_0_elements(62) <= In_wrap_daemon_CP_0_elements(60);
    -- CP-element group 63:  transition  input  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63:  members (6) 
      -- CP-element group 63: 	 branch_block_stmt_31/assign_stmt_120/RPIPE_w_in_buf_119_sample_completed_
      -- CP-element group 63: 	 branch_block_stmt_31/assign_stmt_120/RPIPE_w_in_buf_119_update_start_
      -- CP-element group 63: 	 branch_block_stmt_31/assign_stmt_120/RPIPE_w_in_buf_119_Sample/$exit
      -- CP-element group 63: 	 branch_block_stmt_31/assign_stmt_120/RPIPE_w_in_buf_119_Sample/ra
      -- CP-element group 63: 	 branch_block_stmt_31/assign_stmt_120/RPIPE_w_in_buf_119_Update/$entry
      -- CP-element group 63: 	 branch_block_stmt_31/assign_stmt_120/RPIPE_w_in_buf_119_Update/cr
      -- 
    ra_497_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_w_in_buf_119_inst_ack_0, ack => In_wrap_daemon_CP_0_elements(63)); -- 
    cr_501_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_501_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => In_wrap_daemon_CP_0_elements(63), ack => RPIPE_w_in_buf_119_inst_req_1); -- 
    -- CP-element group 64:  transition  input  output  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	65 
    -- CP-element group 64:  members (6) 
      -- CP-element group 64: 	 branch_block_stmt_31/assign_stmt_120/RPIPE_w_in_buf_119_update_completed_
      -- CP-element group 64: 	 branch_block_stmt_31/assign_stmt_120/RPIPE_w_in_buf_119_Update/$exit
      -- CP-element group 64: 	 branch_block_stmt_31/assign_stmt_120/RPIPE_w_in_buf_119_Update/ca
      -- CP-element group 64: 	 branch_block_stmt_31/assign_stmt_120/WPIPE_e_in_buf_118_sample_start_
      -- CP-element group 64: 	 branch_block_stmt_31/assign_stmt_120/WPIPE_e_in_buf_118_Sample/$entry
      -- CP-element group 64: 	 branch_block_stmt_31/assign_stmt_120/WPIPE_e_in_buf_118_Sample/req
      -- 
    ca_502_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_w_in_buf_119_inst_ack_1, ack => In_wrap_daemon_CP_0_elements(64)); -- 
    req_510_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_510_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => In_wrap_daemon_CP_0_elements(64), ack => WPIPE_e_in_buf_118_inst_req_0); -- 
    -- CP-element group 65:  transition  input  output  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	64 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	66 
    -- CP-element group 65:  members (6) 
      -- CP-element group 65: 	 branch_block_stmt_31/assign_stmt_120/WPIPE_e_in_buf_118_sample_completed_
      -- CP-element group 65: 	 branch_block_stmt_31/assign_stmt_120/WPIPE_e_in_buf_118_update_start_
      -- CP-element group 65: 	 branch_block_stmt_31/assign_stmt_120/WPIPE_e_in_buf_118_Sample/$exit
      -- CP-element group 65: 	 branch_block_stmt_31/assign_stmt_120/WPIPE_e_in_buf_118_Sample/ack
      -- CP-element group 65: 	 branch_block_stmt_31/assign_stmt_120/WPIPE_e_in_buf_118_Update/$entry
      -- CP-element group 65: 	 branch_block_stmt_31/assign_stmt_120/WPIPE_e_in_buf_118_Update/req
      -- 
    ack_511_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_e_in_buf_118_inst_ack_0, ack => In_wrap_daemon_CP_0_elements(65)); -- 
    req_515_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_515_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => In_wrap_daemon_CP_0_elements(65), ack => WPIPE_e_in_buf_118_inst_req_1); -- 
    -- CP-element group 66:  transition  input  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	65 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	61 
    -- CP-element group 66:  members (4) 
      -- CP-element group 66: 	 branch_block_stmt_31/assign_stmt_120/$exit
      -- CP-element group 66: 	 branch_block_stmt_31/assign_stmt_120/WPIPE_e_in_buf_118_update_completed_
      -- CP-element group 66: 	 branch_block_stmt_31/assign_stmt_120/WPIPE_e_in_buf_118_Update/$exit
      -- CP-element group 66: 	 branch_block_stmt_31/assign_stmt_120/WPIPE_e_in_buf_118_Update/ack
      -- 
    ack_516_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_e_in_buf_118_inst_ack_1, ack => In_wrap_daemon_CP_0_elements(66)); -- 
    -- CP-element group 67:  place  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	59 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	69 
    -- CP-element group 67:  members (1) 
      -- CP-element group 67: 	 branch_block_stmt_31/assign_stmt_124__entry__
      -- 
    In_wrap_daemon_CP_0_elements(67) <= In_wrap_daemon_CP_0_elements(59);
    -- CP-element group 68:  place  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	73 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	10 
    -- CP-element group 68:  members (1) 
      -- CP-element group 68: 	 branch_block_stmt_31/assign_stmt_124__exit__
      -- 
    In_wrap_daemon_CP_0_elements(68) <= In_wrap_daemon_CP_0_elements(73);
    -- CP-element group 69:  transition  output  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	67 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	70 
    -- CP-element group 69:  members (4) 
      -- CP-element group 69: 	 branch_block_stmt_31/assign_stmt_124/$entry
      -- CP-element group 69: 	 branch_block_stmt_31/assign_stmt_124/RPIPE_w_in_buf_123_sample_start_
      -- CP-element group 69: 	 branch_block_stmt_31/assign_stmt_124/RPIPE_w_in_buf_123_Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_31/assign_stmt_124/RPIPE_w_in_buf_123_Sample/rr
      -- 
    rr_529_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_529_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => In_wrap_daemon_CP_0_elements(69), ack => RPIPE_w_in_buf_123_inst_req_0); -- 
    In_wrap_daemon_CP_0_elements(69) <= In_wrap_daemon_CP_0_elements(67);
    -- CP-element group 70:  transition  input  output  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	69 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70:  members (6) 
      -- CP-element group 70: 	 branch_block_stmt_31/assign_stmt_124/RPIPE_w_in_buf_123_sample_completed_
      -- CP-element group 70: 	 branch_block_stmt_31/assign_stmt_124/RPIPE_w_in_buf_123_update_start_
      -- CP-element group 70: 	 branch_block_stmt_31/assign_stmt_124/RPIPE_w_in_buf_123_Sample/$exit
      -- CP-element group 70: 	 branch_block_stmt_31/assign_stmt_124/RPIPE_w_in_buf_123_Sample/ra
      -- CP-element group 70: 	 branch_block_stmt_31/assign_stmt_124/RPIPE_w_in_buf_123_Update/$entry
      -- CP-element group 70: 	 branch_block_stmt_31/assign_stmt_124/RPIPE_w_in_buf_123_Update/cr
      -- 
    ra_530_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_w_in_buf_123_inst_ack_0, ack => In_wrap_daemon_CP_0_elements(70)); -- 
    cr_534_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_534_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => In_wrap_daemon_CP_0_elements(70), ack => RPIPE_w_in_buf_123_inst_req_1); -- 
    -- CP-element group 71:  transition  input  output  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	72 
    -- CP-element group 71:  members (6) 
      -- CP-element group 71: 	 branch_block_stmt_31/assign_stmt_124/RPIPE_w_in_buf_123_update_completed_
      -- CP-element group 71: 	 branch_block_stmt_31/assign_stmt_124/RPIPE_w_in_buf_123_Update/$exit
      -- CP-element group 71: 	 branch_block_stmt_31/assign_stmt_124/RPIPE_w_in_buf_123_Update/ca
      -- CP-element group 71: 	 branch_block_stmt_31/assign_stmt_124/WPIPE_d_in_buf_122_sample_start_
      -- CP-element group 71: 	 branch_block_stmt_31/assign_stmt_124/WPIPE_d_in_buf_122_Sample/$entry
      -- CP-element group 71: 	 branch_block_stmt_31/assign_stmt_124/WPIPE_d_in_buf_122_Sample/req
      -- 
    ca_535_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_w_in_buf_123_inst_ack_1, ack => In_wrap_daemon_CP_0_elements(71)); -- 
    req_543_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_543_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => In_wrap_daemon_CP_0_elements(71), ack => WPIPE_d_in_buf_122_inst_req_0); -- 
    -- CP-element group 72:  transition  input  output  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	71 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	73 
    -- CP-element group 72:  members (6) 
      -- CP-element group 72: 	 branch_block_stmt_31/assign_stmt_124/WPIPE_d_in_buf_122_sample_completed_
      -- CP-element group 72: 	 branch_block_stmt_31/assign_stmt_124/WPIPE_d_in_buf_122_update_start_
      -- CP-element group 72: 	 branch_block_stmt_31/assign_stmt_124/WPIPE_d_in_buf_122_Sample/$exit
      -- CP-element group 72: 	 branch_block_stmt_31/assign_stmt_124/WPIPE_d_in_buf_122_Sample/ack
      -- CP-element group 72: 	 branch_block_stmt_31/assign_stmt_124/WPIPE_d_in_buf_122_Update/$entry
      -- CP-element group 72: 	 branch_block_stmt_31/assign_stmt_124/WPIPE_d_in_buf_122_Update/req
      -- 
    ack_544_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_d_in_buf_122_inst_ack_0, ack => In_wrap_daemon_CP_0_elements(72)); -- 
    req_548_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_548_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => In_wrap_daemon_CP_0_elements(72), ack => WPIPE_d_in_buf_122_inst_req_1); -- 
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	72 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	68 
    -- CP-element group 73:  members (4) 
      -- CP-element group 73: 	 branch_block_stmt_31/assign_stmt_124/$exit
      -- CP-element group 73: 	 branch_block_stmt_31/assign_stmt_124/WPIPE_d_in_buf_122_update_completed_
      -- CP-element group 73: 	 branch_block_stmt_31/assign_stmt_124/WPIPE_d_in_buf_122_Update/$exit
      -- CP-element group 73: 	 branch_block_stmt_31/assign_stmt_124/WPIPE_d_in_buf_122_Update/ack
      -- 
    ack_549_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_d_in_buf_122_inst_ack_1, ack => In_wrap_daemon_CP_0_elements(73)); -- 
    -- CP-element group 74:  transition  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	10 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	11 
    -- CP-element group 74:  members (18) 
      -- CP-element group 74: 	 branch_block_stmt_31/assign_stmt_130/$entry
      -- CP-element group 74: 	 branch_block_stmt_31/assign_stmt_130/$exit
      -- CP-element group 74: 	 branch_block_stmt_31/assign_stmt_130/ADD_u15_u15_129_sample_start_
      -- CP-element group 74: 	 branch_block_stmt_31/assign_stmt_130/ADD_u15_u15_129_sample_completed_
      -- CP-element group 74: 	 branch_block_stmt_31/assign_stmt_130/ADD_u15_u15_129_update_start_
      -- CP-element group 74: 	 branch_block_stmt_31/assign_stmt_130/ADD_u15_u15_129_update_completed_
      -- CP-element group 74: 	 branch_block_stmt_31/assign_stmt_130/R_count_var_127_sample_start_
      -- CP-element group 74: 	 branch_block_stmt_31/assign_stmt_130/R_count_var_127_sample_completed_
      -- CP-element group 74: 	 branch_block_stmt_31/assign_stmt_130/R_count_var_127_update_start_
      -- CP-element group 74: 	 branch_block_stmt_31/assign_stmt_130/R_count_var_127_update_completed_
      -- CP-element group 74: 	 branch_block_stmt_31/assign_stmt_130/ADD_u15_u15_129_Sample/$entry
      -- CP-element group 74: 	 branch_block_stmt_31/assign_stmt_130/ADD_u15_u15_129_Sample/$exit
      -- CP-element group 74: 	 branch_block_stmt_31/assign_stmt_130/ADD_u15_u15_129_Sample/rr
      -- CP-element group 74: 	 branch_block_stmt_31/assign_stmt_130/ADD_u15_u15_129_Sample/ra
      -- CP-element group 74: 	 branch_block_stmt_31/assign_stmt_130/ADD_u15_u15_129_Update/$entry
      -- CP-element group 74: 	 branch_block_stmt_31/assign_stmt_130/ADD_u15_u15_129_Update/$exit
      -- CP-element group 74: 	 branch_block_stmt_31/assign_stmt_130/ADD_u15_u15_129_Update/cr
      -- CP-element group 74: 	 branch_block_stmt_31/assign_stmt_130/ADD_u15_u15_129_Update/ca
      -- 
    In_wrap_daemon_CP_0_elements(74) <= In_wrap_daemon_CP_0_elements(10);
    -- CP-element group 75:  transition  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	11 
    -- CP-element group 75: successors 
    -- CP-element group 75:  members (1) 
      -- CP-element group 75: 	 branch_block_stmt_31/if_stmt_131_dead_link/$entry
      -- 
    In_wrap_daemon_CP_0_elements(75) <= In_wrap_daemon_CP_0_elements(11);
    -- CP-element group 76:  transition  output  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	11 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	77 
    -- CP-element group 76:  members (17) 
      -- CP-element group 76: 	 branch_block_stmt_31/if_stmt_131_eval_test/$entry
      -- CP-element group 76: 	 branch_block_stmt_31/if_stmt_131_eval_test/$exit
      -- CP-element group 76: 	 branch_block_stmt_31/if_stmt_131_eval_test/ULT_u15_u1_134/$entry
      -- CP-element group 76: 	 branch_block_stmt_31/if_stmt_131_eval_test/ULT_u15_u1_134/$exit
      -- CP-element group 76: 	 branch_block_stmt_31/if_stmt_131_eval_test/ULT_u15_u1_134/ULT_u15_u1_134_inputs/$entry
      -- CP-element group 76: 	 branch_block_stmt_31/if_stmt_131_eval_test/ULT_u15_u1_134/ULT_u15_u1_134_inputs/$exit
      -- CP-element group 76: 	 branch_block_stmt_31/if_stmt_131_eval_test/ULT_u15_u1_134/SplitProtocol/$entry
      -- CP-element group 76: 	 branch_block_stmt_31/if_stmt_131_eval_test/ULT_u15_u1_134/SplitProtocol/$exit
      -- CP-element group 76: 	 branch_block_stmt_31/if_stmt_131_eval_test/ULT_u15_u1_134/SplitProtocol/Sample/$entry
      -- CP-element group 76: 	 branch_block_stmt_31/if_stmt_131_eval_test/ULT_u15_u1_134/SplitProtocol/Sample/$exit
      -- CP-element group 76: 	 branch_block_stmt_31/if_stmt_131_eval_test/ULT_u15_u1_134/SplitProtocol/Sample/rr
      -- CP-element group 76: 	 branch_block_stmt_31/if_stmt_131_eval_test/ULT_u15_u1_134/SplitProtocol/Sample/ra
      -- CP-element group 76: 	 branch_block_stmt_31/if_stmt_131_eval_test/ULT_u15_u1_134/SplitProtocol/Update/$entry
      -- CP-element group 76: 	 branch_block_stmt_31/if_stmt_131_eval_test/ULT_u15_u1_134/SplitProtocol/Update/$exit
      -- CP-element group 76: 	 branch_block_stmt_31/if_stmt_131_eval_test/ULT_u15_u1_134/SplitProtocol/Update/cr
      -- CP-element group 76: 	 branch_block_stmt_31/if_stmt_131_eval_test/ULT_u15_u1_134/SplitProtocol/Update/ca
      -- CP-element group 76: 	 branch_block_stmt_31/if_stmt_131_eval_test/branch_req
      -- 
    branch_req_597_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_597_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => In_wrap_daemon_CP_0_elements(76), ack => if_stmt_131_branch_req_0); -- 
    In_wrap_daemon_CP_0_elements(76) <= In_wrap_daemon_CP_0_elements(11);
    -- CP-element group 77:  branch  place  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	76 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	78 
    -- CP-element group 77: 	80 
    -- CP-element group 77:  members (1) 
      -- CP-element group 77: 	 branch_block_stmt_31/ULT_u15_u1_134_place
      -- 
    In_wrap_daemon_CP_0_elements(77) <= In_wrap_daemon_CP_0_elements(76);
    -- CP-element group 78:  transition  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	77 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	79 
    -- CP-element group 78:  members (1) 
      -- CP-element group 78: 	 branch_block_stmt_31/if_stmt_131_if_link/$entry
      -- 
    In_wrap_daemon_CP_0_elements(78) <= In_wrap_daemon_CP_0_elements(77);
    -- CP-element group 79:  transition  input  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	78 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	82 
    -- CP-element group 79:  members (2) 
      -- CP-element group 79: 	 branch_block_stmt_31/if_stmt_131_if_link/$exit
      -- CP-element group 79: 	 branch_block_stmt_31/if_stmt_131_if_link/if_choice_transition
      -- 
    if_choice_transition_602_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_131_branch_ack_1, ack => In_wrap_daemon_CP_0_elements(79)); -- 
    -- CP-element group 80:  transition  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	77 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	81 
    -- CP-element group 80:  members (1) 
      -- CP-element group 80: 	 branch_block_stmt_31/if_stmt_131_else_link/$entry
      -- 
    In_wrap_daemon_CP_0_elements(80) <= In_wrap_daemon_CP_0_elements(77);
    -- CP-element group 81:  transition  input  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	80 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	83 
    -- CP-element group 81:  members (2) 
      -- CP-element group 81: 	 branch_block_stmt_31/if_stmt_131_else_link/$exit
      -- CP-element group 81: 	 branch_block_stmt_31/if_stmt_131_else_link/else_choice_transition
      -- 
    else_choice_transition_606_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_131_branch_ack_0, ack => In_wrap_daemon_CP_0_elements(81)); -- 
    -- CP-element group 82:  place  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	79 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	125 
    -- CP-element group 82:  members (1) 
      -- CP-element group 82: 	 branch_block_stmt_31/loop1
      -- 
    In_wrap_daemon_CP_0_elements(82) <= In_wrap_daemon_CP_0_elements(79);
    -- CP-element group 83:  branch  place  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	81 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	85 
    -- CP-element group 83: 	86 
    -- CP-element group 83:  members (1) 
      -- CP-element group 83: 	 branch_block_stmt_31/if_stmt_137__entry__
      -- 
    In_wrap_daemon_CP_0_elements(83) <= In_wrap_daemon_CP_0_elements(81);
    -- CP-element group 84:  merge  place  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	91 
    -- CP-element group 84: 	96 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	132 
    -- CP-element group 84:  members (3) 
      -- CP-element group 84: 	 branch_block_stmt_31/branch_block_stmt_31__exit__
      -- CP-element group 84: 	 branch_block_stmt_31/if_stmt_131__exit__
      -- CP-element group 84: 	 branch_block_stmt_31/if_stmt_137__exit__
      -- 
    In_wrap_daemon_CP_0_elements(84) <= OrReduce(In_wrap_daemon_CP_0_elements(91) & In_wrap_daemon_CP_0_elements(96));
    -- CP-element group 85:  transition  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	83 
    -- CP-element group 85: successors 
    -- CP-element group 85:  members (1) 
      -- CP-element group 85: 	 branch_block_stmt_31/if_stmt_137_dead_link/$entry
      -- 
    In_wrap_daemon_CP_0_elements(85) <= In_wrap_daemon_CP_0_elements(83);
    -- CP-element group 86:  transition  output  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	83 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	87 
    -- CP-element group 86:  members (17) 
      -- CP-element group 86: 	 branch_block_stmt_31/if_stmt_137_eval_test/$entry
      -- CP-element group 86: 	 branch_block_stmt_31/if_stmt_137_eval_test/$exit
      -- CP-element group 86: 	 branch_block_stmt_31/if_stmt_137_eval_test/ULT_u15_u1_140/$entry
      -- CP-element group 86: 	 branch_block_stmt_31/if_stmt_137_eval_test/ULT_u15_u1_140/$exit
      -- CP-element group 86: 	 branch_block_stmt_31/if_stmt_137_eval_test/ULT_u15_u1_140/ULT_u15_u1_140_inputs/$entry
      -- CP-element group 86: 	 branch_block_stmt_31/if_stmt_137_eval_test/ULT_u15_u1_140/ULT_u15_u1_140_inputs/$exit
      -- CP-element group 86: 	 branch_block_stmt_31/if_stmt_137_eval_test/ULT_u15_u1_140/SplitProtocol/$entry
      -- CP-element group 86: 	 branch_block_stmt_31/if_stmt_137_eval_test/ULT_u15_u1_140/SplitProtocol/$exit
      -- CP-element group 86: 	 branch_block_stmt_31/if_stmt_137_eval_test/ULT_u15_u1_140/SplitProtocol/Sample/$entry
      -- CP-element group 86: 	 branch_block_stmt_31/if_stmt_137_eval_test/ULT_u15_u1_140/SplitProtocol/Sample/$exit
      -- CP-element group 86: 	 branch_block_stmt_31/if_stmt_137_eval_test/ULT_u15_u1_140/SplitProtocol/Sample/rr
      -- CP-element group 86: 	 branch_block_stmt_31/if_stmt_137_eval_test/ULT_u15_u1_140/SplitProtocol/Sample/ra
      -- CP-element group 86: 	 branch_block_stmt_31/if_stmt_137_eval_test/ULT_u15_u1_140/SplitProtocol/Update/$entry
      -- CP-element group 86: 	 branch_block_stmt_31/if_stmt_137_eval_test/ULT_u15_u1_140/SplitProtocol/Update/$exit
      -- CP-element group 86: 	 branch_block_stmt_31/if_stmt_137_eval_test/ULT_u15_u1_140/SplitProtocol/Update/cr
      -- CP-element group 86: 	 branch_block_stmt_31/if_stmt_137_eval_test/ULT_u15_u1_140/SplitProtocol/Update/ca
      -- CP-element group 86: 	 branch_block_stmt_31/if_stmt_137_eval_test/branch_req
      -- 
    branch_req_636_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_636_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => In_wrap_daemon_CP_0_elements(86), ack => if_stmt_137_branch_req_0); -- 
    In_wrap_daemon_CP_0_elements(86) <= In_wrap_daemon_CP_0_elements(83);
    -- CP-element group 87:  branch  place  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	86 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87: 	90 
    -- CP-element group 87:  members (1) 
      -- CP-element group 87: 	 branch_block_stmt_31/ULT_u15_u1_140_place
      -- 
    In_wrap_daemon_CP_0_elements(87) <= In_wrap_daemon_CP_0_elements(86);
    -- CP-element group 88:  transition  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	87 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	89 
    -- CP-element group 88:  members (1) 
      -- CP-element group 88: 	 branch_block_stmt_31/if_stmt_137_if_link/$entry
      -- 
    In_wrap_daemon_CP_0_elements(88) <= In_wrap_daemon_CP_0_elements(87);
    -- CP-element group 89:  transition  input  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	88 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	92 
    -- CP-element group 89:  members (2) 
      -- CP-element group 89: 	 branch_block_stmt_31/if_stmt_137_if_link/$exit
      -- CP-element group 89: 	 branch_block_stmt_31/if_stmt_137_if_link/if_choice_transition
      -- 
    if_choice_transition_641_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_137_branch_ack_1, ack => In_wrap_daemon_CP_0_elements(89)); -- 
    -- CP-element group 90:  transition  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	87 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	91 
    -- CP-element group 90:  members (1) 
      -- CP-element group 90: 	 branch_block_stmt_31/if_stmt_137_else_link/$entry
      -- 
    In_wrap_daemon_CP_0_elements(90) <= In_wrap_daemon_CP_0_elements(87);
    -- CP-element group 91:  transition  input  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	90 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	84 
    -- CP-element group 91:  members (2) 
      -- CP-element group 91: 	 branch_block_stmt_31/if_stmt_137_else_link/$exit
      -- CP-element group 91: 	 branch_block_stmt_31/if_stmt_137_else_link/else_choice_transition
      -- 
    else_choice_transition_645_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_137_branch_ack_0, ack => In_wrap_daemon_CP_0_elements(91)); -- 
    -- CP-element group 92:  branch  place  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	89 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	111 
    -- CP-element group 92: 	112 
    -- CP-element group 92:  members (1) 
      -- CP-element group 92: 	 branch_block_stmt_31/merge_stmt_141__entry__
      -- 
    In_wrap_daemon_CP_0_elements(92) <= In_wrap_daemon_CP_0_elements(89);
    -- CP-element group 93:  merge  place  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	122 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	97 
    -- CP-element group 93:  members (2) 
      -- CP-element group 93: 	 branch_block_stmt_31/merge_stmt_141__exit__
      -- CP-element group 93: 	 branch_block_stmt_31/assign_stmt_149__entry__
      -- 
    In_wrap_daemon_CP_0_elements(93) <= In_wrap_daemon_CP_0_elements(122);
    -- CP-element group 94:  place  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	101 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	102 
    -- CP-element group 94:  members (2) 
      -- CP-element group 94: 	 branch_block_stmt_31/assign_stmt_149__exit__
      -- CP-element group 94: 	 branch_block_stmt_31/assign_stmt_154__entry__
      -- 
    In_wrap_daemon_CP_0_elements(94) <= In_wrap_daemon_CP_0_elements(101);
    -- CP-element group 95:  branch  place  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	102 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	103 
    -- CP-element group 95: 	104 
    -- CP-element group 95:  members (2) 
      -- CP-element group 95: 	 branch_block_stmt_31/assign_stmt_154__exit__
      -- CP-element group 95: 	 branch_block_stmt_31/if_stmt_155__entry__
      -- 
    In_wrap_daemon_CP_0_elements(95) <= In_wrap_daemon_CP_0_elements(102);
    -- CP-element group 96:  merge  place  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	109 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	84 
    -- CP-element group 96:  members (1) 
      -- CP-element group 96: 	 branch_block_stmt_31/if_stmt_155__exit__
      -- 
    In_wrap_daemon_CP_0_elements(96) <= In_wrap_daemon_CP_0_elements(109);
    -- CP-element group 97:  transition  output  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	93 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	98 
    -- CP-element group 97:  members (4) 
      -- CP-element group 97: 	 branch_block_stmt_31/assign_stmt_149/$entry
      -- CP-element group 97: 	 branch_block_stmt_31/assign_stmt_149/RPIPE_w_in_buf_148_sample_start_
      -- CP-element group 97: 	 branch_block_stmt_31/assign_stmt_149/RPIPE_w_in_buf_148_Sample/$entry
      -- CP-element group 97: 	 branch_block_stmt_31/assign_stmt_149/RPIPE_w_in_buf_148_Sample/rr
      -- 
    rr_664_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_664_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => In_wrap_daemon_CP_0_elements(97), ack => RPIPE_w_in_buf_148_inst_req_0); -- 
    In_wrap_daemon_CP_0_elements(97) <= In_wrap_daemon_CP_0_elements(93);
    -- CP-element group 98:  transition  input  output  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	97 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	99 
    -- CP-element group 98:  members (6) 
      -- CP-element group 98: 	 branch_block_stmt_31/assign_stmt_149/RPIPE_w_in_buf_148_sample_completed_
      -- CP-element group 98: 	 branch_block_stmt_31/assign_stmt_149/RPIPE_w_in_buf_148_update_start_
      -- CP-element group 98: 	 branch_block_stmt_31/assign_stmt_149/RPIPE_w_in_buf_148_Sample/$exit
      -- CP-element group 98: 	 branch_block_stmt_31/assign_stmt_149/RPIPE_w_in_buf_148_Sample/ra
      -- CP-element group 98: 	 branch_block_stmt_31/assign_stmt_149/RPIPE_w_in_buf_148_Update/$entry
      -- CP-element group 98: 	 branch_block_stmt_31/assign_stmt_149/RPIPE_w_in_buf_148_Update/cr
      -- 
    ra_665_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_w_in_buf_148_inst_ack_0, ack => In_wrap_daemon_CP_0_elements(98)); -- 
    cr_669_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_669_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => In_wrap_daemon_CP_0_elements(98), ack => RPIPE_w_in_buf_148_inst_req_1); -- 
    -- CP-element group 99:  transition  input  output  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	98 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	100 
    -- CP-element group 99:  members (6) 
      -- CP-element group 99: 	 branch_block_stmt_31/assign_stmt_149/RPIPE_w_in_buf_148_update_completed_
      -- CP-element group 99: 	 branch_block_stmt_31/assign_stmt_149/RPIPE_w_in_buf_148_Update/$exit
      -- CP-element group 99: 	 branch_block_stmt_31/assign_stmt_149/RPIPE_w_in_buf_148_Update/ca
      -- CP-element group 99: 	 branch_block_stmt_31/assign_stmt_149/WPIPE_out_wrap_data_147_sample_start_
      -- CP-element group 99: 	 branch_block_stmt_31/assign_stmt_149/WPIPE_out_wrap_data_147_Sample/$entry
      -- CP-element group 99: 	 branch_block_stmt_31/assign_stmt_149/WPIPE_out_wrap_data_147_Sample/req
      -- 
    ca_670_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_w_in_buf_148_inst_ack_1, ack => In_wrap_daemon_CP_0_elements(99)); -- 
    req_678_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_678_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => In_wrap_daemon_CP_0_elements(99), ack => WPIPE_out_wrap_data_147_inst_req_0); -- 
    -- CP-element group 100:  transition  input  output  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	99 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	101 
    -- CP-element group 100:  members (6) 
      -- CP-element group 100: 	 branch_block_stmt_31/assign_stmt_149/WPIPE_out_wrap_data_147_sample_completed_
      -- CP-element group 100: 	 branch_block_stmt_31/assign_stmt_149/WPIPE_out_wrap_data_147_update_start_
      -- CP-element group 100: 	 branch_block_stmt_31/assign_stmt_149/WPIPE_out_wrap_data_147_Sample/$exit
      -- CP-element group 100: 	 branch_block_stmt_31/assign_stmt_149/WPIPE_out_wrap_data_147_Sample/ack
      -- CP-element group 100: 	 branch_block_stmt_31/assign_stmt_149/WPIPE_out_wrap_data_147_Update/$entry
      -- CP-element group 100: 	 branch_block_stmt_31/assign_stmt_149/WPIPE_out_wrap_data_147_Update/req
      -- 
    ack_679_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_out_wrap_data_147_inst_ack_0, ack => In_wrap_daemon_CP_0_elements(100)); -- 
    req_683_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_683_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => In_wrap_daemon_CP_0_elements(100), ack => WPIPE_out_wrap_data_147_inst_req_1); -- 
    -- CP-element group 101:  transition  input  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	100 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	94 
    -- CP-element group 101:  members (4) 
      -- CP-element group 101: 	 branch_block_stmt_31/assign_stmt_149/$exit
      -- CP-element group 101: 	 branch_block_stmt_31/assign_stmt_149/WPIPE_out_wrap_data_147_update_completed_
      -- CP-element group 101: 	 branch_block_stmt_31/assign_stmt_149/WPIPE_out_wrap_data_147_Update/$exit
      -- CP-element group 101: 	 branch_block_stmt_31/assign_stmt_149/WPIPE_out_wrap_data_147_Update/ack
      -- 
    ack_684_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_out_wrap_data_147_inst_ack_1, ack => In_wrap_daemon_CP_0_elements(101)); -- 
    -- CP-element group 102:  transition  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	94 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	95 
    -- CP-element group 102:  members (18) 
      -- CP-element group 102: 	 branch_block_stmt_31/assign_stmt_154/$entry
      -- CP-element group 102: 	 branch_block_stmt_31/assign_stmt_154/$exit
      -- CP-element group 102: 	 branch_block_stmt_31/assign_stmt_154/ADD_u15_u15_153_sample_start_
      -- CP-element group 102: 	 branch_block_stmt_31/assign_stmt_154/ADD_u15_u15_153_sample_completed_
      -- CP-element group 102: 	 branch_block_stmt_31/assign_stmt_154/ADD_u15_u15_153_update_start_
      -- CP-element group 102: 	 branch_block_stmt_31/assign_stmt_154/ADD_u15_u15_153_update_completed_
      -- CP-element group 102: 	 branch_block_stmt_31/assign_stmt_154/R_count_var2_151_sample_start_
      -- CP-element group 102: 	 branch_block_stmt_31/assign_stmt_154/R_count_var2_151_sample_completed_
      -- CP-element group 102: 	 branch_block_stmt_31/assign_stmt_154/R_count_var2_151_update_start_
      -- CP-element group 102: 	 branch_block_stmt_31/assign_stmt_154/R_count_var2_151_update_completed_
      -- CP-element group 102: 	 branch_block_stmt_31/assign_stmt_154/ADD_u15_u15_153_Sample/$entry
      -- CP-element group 102: 	 branch_block_stmt_31/assign_stmt_154/ADD_u15_u15_153_Sample/$exit
      -- CP-element group 102: 	 branch_block_stmt_31/assign_stmt_154/ADD_u15_u15_153_Sample/rr
      -- CP-element group 102: 	 branch_block_stmt_31/assign_stmt_154/ADD_u15_u15_153_Sample/ra
      -- CP-element group 102: 	 branch_block_stmt_31/assign_stmt_154/ADD_u15_u15_153_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_31/assign_stmt_154/ADD_u15_u15_153_Update/$exit
      -- CP-element group 102: 	 branch_block_stmt_31/assign_stmt_154/ADD_u15_u15_153_Update/cr
      -- CP-element group 102: 	 branch_block_stmt_31/assign_stmt_154/ADD_u15_u15_153_Update/ca
      -- 
    In_wrap_daemon_CP_0_elements(102) <= In_wrap_daemon_CP_0_elements(94);
    -- CP-element group 103:  transition  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	95 
    -- CP-element group 103: successors 
    -- CP-element group 103:  members (1) 
      -- CP-element group 103: 	 branch_block_stmt_31/if_stmt_155_dead_link/$entry
      -- 
    In_wrap_daemon_CP_0_elements(103) <= In_wrap_daemon_CP_0_elements(95);
    -- CP-element group 104:  transition  output  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	95 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	105 
    -- CP-element group 104:  members (17) 
      -- CP-element group 104: 	 branch_block_stmt_31/if_stmt_155_eval_test/$entry
      -- CP-element group 104: 	 branch_block_stmt_31/if_stmt_155_eval_test/$exit
      -- CP-element group 104: 	 branch_block_stmt_31/if_stmt_155_eval_test/ULT_u15_u1_158/$entry
      -- CP-element group 104: 	 branch_block_stmt_31/if_stmt_155_eval_test/ULT_u15_u1_158/$exit
      -- CP-element group 104: 	 branch_block_stmt_31/if_stmt_155_eval_test/ULT_u15_u1_158/ULT_u15_u1_158_inputs/$entry
      -- CP-element group 104: 	 branch_block_stmt_31/if_stmt_155_eval_test/ULT_u15_u1_158/ULT_u15_u1_158_inputs/$exit
      -- CP-element group 104: 	 branch_block_stmt_31/if_stmt_155_eval_test/ULT_u15_u1_158/SplitProtocol/$entry
      -- CP-element group 104: 	 branch_block_stmt_31/if_stmt_155_eval_test/ULT_u15_u1_158/SplitProtocol/$exit
      -- CP-element group 104: 	 branch_block_stmt_31/if_stmt_155_eval_test/ULT_u15_u1_158/SplitProtocol/Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_31/if_stmt_155_eval_test/ULT_u15_u1_158/SplitProtocol/Sample/$exit
      -- CP-element group 104: 	 branch_block_stmt_31/if_stmt_155_eval_test/ULT_u15_u1_158/SplitProtocol/Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_31/if_stmt_155_eval_test/ULT_u15_u1_158/SplitProtocol/Sample/ra
      -- CP-element group 104: 	 branch_block_stmt_31/if_stmt_155_eval_test/ULT_u15_u1_158/SplitProtocol/Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_31/if_stmt_155_eval_test/ULT_u15_u1_158/SplitProtocol/Update/$exit
      -- CP-element group 104: 	 branch_block_stmt_31/if_stmt_155_eval_test/ULT_u15_u1_158/SplitProtocol/Update/cr
      -- CP-element group 104: 	 branch_block_stmt_31/if_stmt_155_eval_test/ULT_u15_u1_158/SplitProtocol/Update/ca
      -- CP-element group 104: 	 branch_block_stmt_31/if_stmt_155_eval_test/branch_req
      -- 
    branch_req_732_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_732_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => In_wrap_daemon_CP_0_elements(104), ack => if_stmt_155_branch_req_0); -- 
    In_wrap_daemon_CP_0_elements(104) <= In_wrap_daemon_CP_0_elements(95);
    -- CP-element group 105:  branch  place  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	104 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	106 
    -- CP-element group 105: 	108 
    -- CP-element group 105:  members (1) 
      -- CP-element group 105: 	 branch_block_stmt_31/ULT_u15_u1_158_place
      -- 
    In_wrap_daemon_CP_0_elements(105) <= In_wrap_daemon_CP_0_elements(104);
    -- CP-element group 106:  transition  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	105 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	107 
    -- CP-element group 106:  members (1) 
      -- CP-element group 106: 	 branch_block_stmt_31/if_stmt_155_if_link/$entry
      -- 
    In_wrap_daemon_CP_0_elements(106) <= In_wrap_daemon_CP_0_elements(105);
    -- CP-element group 107:  transition  input  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	106 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	110 
    -- CP-element group 107:  members (2) 
      -- CP-element group 107: 	 branch_block_stmt_31/if_stmt_155_if_link/$exit
      -- CP-element group 107: 	 branch_block_stmt_31/if_stmt_155_if_link/if_choice_transition
      -- 
    if_choice_transition_737_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_155_branch_ack_1, ack => In_wrap_daemon_CP_0_elements(107)); -- 
    -- CP-element group 108:  transition  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	105 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	109 
    -- CP-element group 108:  members (1) 
      -- CP-element group 108: 	 branch_block_stmt_31/if_stmt_155_else_link/$entry
      -- 
    In_wrap_daemon_CP_0_elements(108) <= In_wrap_daemon_CP_0_elements(105);
    -- CP-element group 109:  transition  input  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	108 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	96 
    -- CP-element group 109:  members (2) 
      -- CP-element group 109: 	 branch_block_stmt_31/if_stmt_155_else_link/$exit
      -- CP-element group 109: 	 branch_block_stmt_31/if_stmt_155_else_link/else_choice_transition
      -- 
    else_choice_transition_741_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_155_branch_ack_0, ack => In_wrap_daemon_CP_0_elements(109)); -- 
    -- CP-element group 110:  place  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	107 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	116 
    -- CP-element group 110:  members (1) 
      -- CP-element group 110: 	 branch_block_stmt_31/loop2
      -- 
    In_wrap_daemon_CP_0_elements(110) <= In_wrap_daemon_CP_0_elements(107);
    -- CP-element group 111:  transition  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	92 
    -- CP-element group 111: successors 
    -- CP-element group 111:  members (1) 
      -- CP-element group 111: 	 branch_block_stmt_31/merge_stmt_141_dead_link/$entry
      -- 
    In_wrap_daemon_CP_0_elements(111) <= In_wrap_daemon_CP_0_elements(92);
    -- CP-element group 112:  fork  transition  output  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	92 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	113 
    -- CP-element group 112: 	114 
    -- CP-element group 112:  members (8) 
      -- CP-element group 112: 	 branch_block_stmt_31/merge_stmt_141__entry___PhiReq/$entry
      -- CP-element group 112: 	 branch_block_stmt_31/merge_stmt_141__entry___PhiReq/phi_stmt_142/$entry
      -- CP-element group 112: 	 branch_block_stmt_31/merge_stmt_141__entry___PhiReq/phi_stmt_142/phi_stmt_142_sources/$entry
      -- CP-element group 112: 	 branch_block_stmt_31/merge_stmt_141__entry___PhiReq/phi_stmt_142/phi_stmt_142_sources/Interlock/$entry
      -- CP-element group 112: 	 branch_block_stmt_31/merge_stmt_141__entry___PhiReq/phi_stmt_142/phi_stmt_142_sources/Interlock/Sample/$entry
      -- CP-element group 112: 	 branch_block_stmt_31/merge_stmt_141__entry___PhiReq/phi_stmt_142/phi_stmt_142_sources/Interlock/Sample/req
      -- CP-element group 112: 	 branch_block_stmt_31/merge_stmt_141__entry___PhiReq/phi_stmt_142/phi_stmt_142_sources/Interlock/Update/$entry
      -- CP-element group 112: 	 branch_block_stmt_31/merge_stmt_141__entry___PhiReq/phi_stmt_142/phi_stmt_142_sources/Interlock/Update/req
      -- 
    req_762_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_762_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => In_wrap_daemon_CP_0_elements(112), ack => n_count_var_130_144_buf_req_0); -- 
    req_767_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_767_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => In_wrap_daemon_CP_0_elements(112), ack => n_count_var_130_144_buf_req_1); -- 
    In_wrap_daemon_CP_0_elements(112) <= In_wrap_daemon_CP_0_elements(92);
    -- CP-element group 113:  transition  input  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	112 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	115 
    -- CP-element group 113:  members (2) 
      -- CP-element group 113: 	 branch_block_stmt_31/merge_stmt_141__entry___PhiReq/phi_stmt_142/phi_stmt_142_sources/Interlock/Sample/$exit
      -- CP-element group 113: 	 branch_block_stmt_31/merge_stmt_141__entry___PhiReq/phi_stmt_142/phi_stmt_142_sources/Interlock/Sample/ack
      -- 
    ack_763_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_count_var_130_144_buf_ack_0, ack => In_wrap_daemon_CP_0_elements(113)); -- 
    -- CP-element group 114:  transition  input  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	112 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	115 
    -- CP-element group 114:  members (2) 
      -- CP-element group 114: 	 branch_block_stmt_31/merge_stmt_141__entry___PhiReq/phi_stmt_142/phi_stmt_142_sources/Interlock/Update/$exit
      -- CP-element group 114: 	 branch_block_stmt_31/merge_stmt_141__entry___PhiReq/phi_stmt_142/phi_stmt_142_sources/Interlock/Update/ack
      -- 
    ack_768_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_count_var_130_144_buf_ack_1, ack => In_wrap_daemon_CP_0_elements(114)); -- 
    -- CP-element group 115:  join  transition  output  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	113 
    -- CP-element group 115: 	114 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	120 
    -- CP-element group 115:  members (5) 
      -- CP-element group 115: 	 branch_block_stmt_31/merge_stmt_141__entry___PhiReq/$exit
      -- CP-element group 115: 	 branch_block_stmt_31/merge_stmt_141__entry___PhiReq/phi_stmt_142/$exit
      -- CP-element group 115: 	 branch_block_stmt_31/merge_stmt_141__entry___PhiReq/phi_stmt_142/phi_stmt_142_sources/$exit
      -- CP-element group 115: 	 branch_block_stmt_31/merge_stmt_141__entry___PhiReq/phi_stmt_142/phi_stmt_142_sources/Interlock/$exit
      -- CP-element group 115: 	 branch_block_stmt_31/merge_stmt_141__entry___PhiReq/phi_stmt_142/phi_stmt_142_req
      -- 
    phi_stmt_142_req_769_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_142_req_769_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => In_wrap_daemon_CP_0_elements(115), ack => phi_stmt_142_req_0); -- 
    In_wrap_daemon_cp_element_group_115: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "In_wrap_daemon_cp_element_group_115"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= In_wrap_daemon_CP_0_elements(113) & In_wrap_daemon_CP_0_elements(114);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => In_wrap_daemon_CP_0_elements(115), clk => clk, reset => reset); --
    end block;
    -- CP-element group 116:  fork  transition  output  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	110 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	117 
    -- CP-element group 116: 	118 
    -- CP-element group 116:  members (8) 
      -- CP-element group 116: 	 branch_block_stmt_31/loop2_PhiReq/phi_stmt_142/phi_stmt_142_sources/Interlock/Update/$entry
      -- CP-element group 116: 	 branch_block_stmt_31/loop2_PhiReq/phi_stmt_142/phi_stmt_142_sources/Interlock/Update/req
      -- CP-element group 116: 	 branch_block_stmt_31/loop2_PhiReq/$entry
      -- CP-element group 116: 	 branch_block_stmt_31/loop2_PhiReq/phi_stmt_142/$entry
      -- CP-element group 116: 	 branch_block_stmt_31/loop2_PhiReq/phi_stmt_142/phi_stmt_142_sources/$entry
      -- CP-element group 116: 	 branch_block_stmt_31/loop2_PhiReq/phi_stmt_142/phi_stmt_142_sources/Interlock/$entry
      -- CP-element group 116: 	 branch_block_stmt_31/loop2_PhiReq/phi_stmt_142/phi_stmt_142_sources/Interlock/Sample/$entry
      -- CP-element group 116: 	 branch_block_stmt_31/loop2_PhiReq/phi_stmt_142/phi_stmt_142_sources/Interlock/Sample/req
      -- 
    req_785_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_785_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => In_wrap_daemon_CP_0_elements(116), ack => n_count_var2_154_145_buf_req_0); -- 
    req_790_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_790_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => In_wrap_daemon_CP_0_elements(116), ack => n_count_var2_154_145_buf_req_1); -- 
    In_wrap_daemon_CP_0_elements(116) <= In_wrap_daemon_CP_0_elements(110);
    -- CP-element group 117:  transition  input  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	116 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	119 
    -- CP-element group 117:  members (2) 
      -- CP-element group 117: 	 branch_block_stmt_31/loop2_PhiReq/phi_stmt_142/phi_stmt_142_sources/Interlock/Sample/$exit
      -- CP-element group 117: 	 branch_block_stmt_31/loop2_PhiReq/phi_stmt_142/phi_stmt_142_sources/Interlock/Sample/ack
      -- 
    ack_786_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_count_var2_154_145_buf_ack_0, ack => In_wrap_daemon_CP_0_elements(117)); -- 
    -- CP-element group 118:  transition  input  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	116 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	119 
    -- CP-element group 118:  members (2) 
      -- CP-element group 118: 	 branch_block_stmt_31/loop2_PhiReq/phi_stmt_142/phi_stmt_142_sources/Interlock/Update/$exit
      -- CP-element group 118: 	 branch_block_stmt_31/loop2_PhiReq/phi_stmt_142/phi_stmt_142_sources/Interlock/Update/ack
      -- 
    ack_791_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 118_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_count_var2_154_145_buf_ack_1, ack => In_wrap_daemon_CP_0_elements(118)); -- 
    -- CP-element group 119:  join  transition  output  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	117 
    -- CP-element group 119: 	118 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	120 
    -- CP-element group 119:  members (5) 
      -- CP-element group 119: 	 branch_block_stmt_31/loop2_PhiReq/phi_stmt_142/phi_stmt_142_req
      -- CP-element group 119: 	 branch_block_stmt_31/loop2_PhiReq/$exit
      -- CP-element group 119: 	 branch_block_stmt_31/loop2_PhiReq/phi_stmt_142/$exit
      -- CP-element group 119: 	 branch_block_stmt_31/loop2_PhiReq/phi_stmt_142/phi_stmt_142_sources/$exit
      -- CP-element group 119: 	 branch_block_stmt_31/loop2_PhiReq/phi_stmt_142/phi_stmt_142_sources/Interlock/$exit
      -- 
    phi_stmt_142_req_792_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_142_req_792_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => In_wrap_daemon_CP_0_elements(119), ack => phi_stmt_142_req_1); -- 
    In_wrap_daemon_cp_element_group_119: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "In_wrap_daemon_cp_element_group_119"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= In_wrap_daemon_CP_0_elements(117) & In_wrap_daemon_CP_0_elements(118);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => In_wrap_daemon_CP_0_elements(119), clk => clk, reset => reset); --
    end block;
    -- CP-element group 120:  merge  place  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	115 
    -- CP-element group 120: 	119 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	121 
    -- CP-element group 120:  members (1) 
      -- CP-element group 120: 	 branch_block_stmt_31/merge_stmt_141_PhiReqMerge
      -- 
    In_wrap_daemon_CP_0_elements(120) <= OrReduce(In_wrap_daemon_CP_0_elements(115) & In_wrap_daemon_CP_0_elements(119));
    -- CP-element group 121:  transition  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	120 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	122 
    -- CP-element group 121:  members (1) 
      -- CP-element group 121: 	 branch_block_stmt_31/merge_stmt_141_PhiAck/$entry
      -- 
    In_wrap_daemon_CP_0_elements(121) <= In_wrap_daemon_CP_0_elements(120);
    -- CP-element group 122:  transition  input  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	121 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	93 
    -- CP-element group 122:  members (2) 
      -- CP-element group 122: 	 branch_block_stmt_31/merge_stmt_141_PhiAck/$exit
      -- CP-element group 122: 	 branch_block_stmt_31/merge_stmt_141_PhiAck/phi_stmt_142_ack
      -- 
    phi_stmt_142_ack_797_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_142_ack_0, ack => In_wrap_daemon_CP_0_elements(122)); -- 
    -- CP-element group 123:  transition  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	8 
    -- CP-element group 123: successors 
    -- CP-element group 123:  members (1) 
      -- CP-element group 123: 	 branch_block_stmt_31/merge_stmt_108_dead_link/$entry
      -- 
    In_wrap_daemon_CP_0_elements(123) <= In_wrap_daemon_CP_0_elements(8);
    -- CP-element group 124:  transition  output  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	8 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	129 
    -- CP-element group 124:  members (7) 
      -- CP-element group 124: 	 branch_block_stmt_31/merge_stmt_108__entry___PhiReq/$entry
      -- CP-element group 124: 	 branch_block_stmt_31/merge_stmt_108__entry___PhiReq/$exit
      -- CP-element group 124: 	 branch_block_stmt_31/merge_stmt_108__entry___PhiReq/phi_stmt_109/$entry
      -- CP-element group 124: 	 branch_block_stmt_31/merge_stmt_108__entry___PhiReq/phi_stmt_109/$exit
      -- CP-element group 124: 	 branch_block_stmt_31/merge_stmt_108__entry___PhiReq/phi_stmt_109/phi_stmt_109_sources/$entry
      -- CP-element group 124: 	 branch_block_stmt_31/merge_stmt_108__entry___PhiReq/phi_stmt_109/phi_stmt_109_sources/$exit
      -- CP-element group 124: 	 branch_block_stmt_31/merge_stmt_108__entry___PhiReq/phi_stmt_109/phi_stmt_109_req
      -- 
    phi_stmt_109_req_811_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_109_req_811_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => In_wrap_daemon_CP_0_elements(124), ack => phi_stmt_109_req_0); -- 
    In_wrap_daemon_CP_0_elements(124) <= In_wrap_daemon_CP_0_elements(8);
    -- CP-element group 125:  fork  transition  output  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	82 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	126 
    -- CP-element group 125: 	127 
    -- CP-element group 125:  members (8) 
      -- CP-element group 125: 	 branch_block_stmt_31/loop1_PhiReq/$entry
      -- CP-element group 125: 	 branch_block_stmt_31/loop1_PhiReq/phi_stmt_109/$entry
      -- CP-element group 125: 	 branch_block_stmt_31/loop1_PhiReq/phi_stmt_109/phi_stmt_109_sources/$entry
      -- CP-element group 125: 	 branch_block_stmt_31/loop1_PhiReq/phi_stmt_109/phi_stmt_109_sources/Interlock/$entry
      -- CP-element group 125: 	 branch_block_stmt_31/loop1_PhiReq/phi_stmt_109/phi_stmt_109_sources/Interlock/Sample/$entry
      -- CP-element group 125: 	 branch_block_stmt_31/loop1_PhiReq/phi_stmt_109/phi_stmt_109_sources/Interlock/Sample/req
      -- CP-element group 125: 	 branch_block_stmt_31/loop1_PhiReq/phi_stmt_109/phi_stmt_109_sources/Interlock/Update/$entry
      -- CP-element group 125: 	 branch_block_stmt_31/loop1_PhiReq/phi_stmt_109/phi_stmt_109_sources/Interlock/Update/req
      -- 
    req_827_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_827_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => In_wrap_daemon_CP_0_elements(125), ack => n_count_var_130_112_buf_req_0); -- 
    req_832_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_832_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => In_wrap_daemon_CP_0_elements(125), ack => n_count_var_130_112_buf_req_1); -- 
    In_wrap_daemon_CP_0_elements(125) <= In_wrap_daemon_CP_0_elements(82);
    -- CP-element group 126:  transition  input  bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	125 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	128 
    -- CP-element group 126:  members (2) 
      -- CP-element group 126: 	 branch_block_stmt_31/loop1_PhiReq/phi_stmt_109/phi_stmt_109_sources/Interlock/Sample/$exit
      -- CP-element group 126: 	 branch_block_stmt_31/loop1_PhiReq/phi_stmt_109/phi_stmt_109_sources/Interlock/Sample/ack
      -- 
    ack_828_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_count_var_130_112_buf_ack_0, ack => In_wrap_daemon_CP_0_elements(126)); -- 
    -- CP-element group 127:  transition  input  bypass 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	125 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	128 
    -- CP-element group 127:  members (2) 
      -- CP-element group 127: 	 branch_block_stmt_31/loop1_PhiReq/phi_stmt_109/phi_stmt_109_sources/Interlock/Update/$exit
      -- CP-element group 127: 	 branch_block_stmt_31/loop1_PhiReq/phi_stmt_109/phi_stmt_109_sources/Interlock/Update/ack
      -- 
    ack_833_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_count_var_130_112_buf_ack_1, ack => In_wrap_daemon_CP_0_elements(127)); -- 
    -- CP-element group 128:  join  transition  output  bypass 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	126 
    -- CP-element group 128: 	127 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	129 
    -- CP-element group 128:  members (5) 
      -- CP-element group 128: 	 branch_block_stmt_31/loop1_PhiReq/$exit
      -- CP-element group 128: 	 branch_block_stmt_31/loop1_PhiReq/phi_stmt_109/$exit
      -- CP-element group 128: 	 branch_block_stmt_31/loop1_PhiReq/phi_stmt_109/phi_stmt_109_sources/$exit
      -- CP-element group 128: 	 branch_block_stmt_31/loop1_PhiReq/phi_stmt_109/phi_stmt_109_sources/Interlock/$exit
      -- CP-element group 128: 	 branch_block_stmt_31/loop1_PhiReq/phi_stmt_109/phi_stmt_109_req
      -- 
    phi_stmt_109_req_834_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_109_req_834_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => In_wrap_daemon_CP_0_elements(128), ack => phi_stmt_109_req_1); -- 
    In_wrap_daemon_cp_element_group_128: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "In_wrap_daemon_cp_element_group_128"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= In_wrap_daemon_CP_0_elements(126) & In_wrap_daemon_CP_0_elements(127);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => In_wrap_daemon_CP_0_elements(128), clk => clk, reset => reset); --
    end block;
    -- CP-element group 129:  merge  place  bypass 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	124 
    -- CP-element group 129: 	128 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	130 
    -- CP-element group 129:  members (1) 
      -- CP-element group 129: 	 branch_block_stmt_31/merge_stmt_108_PhiReqMerge
      -- 
    In_wrap_daemon_CP_0_elements(129) <= OrReduce(In_wrap_daemon_CP_0_elements(124) & In_wrap_daemon_CP_0_elements(128));
    -- CP-element group 130:  transition  bypass 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	129 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	131 
    -- CP-element group 130:  members (1) 
      -- CP-element group 130: 	 branch_block_stmt_31/merge_stmt_108_PhiAck/$entry
      -- 
    In_wrap_daemon_CP_0_elements(130) <= In_wrap_daemon_CP_0_elements(129);
    -- CP-element group 131:  transition  input  bypass 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	130 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	9 
    -- CP-element group 131:  members (2) 
      -- CP-element group 131: 	 branch_block_stmt_31/merge_stmt_108_PhiAck/$exit
      -- CP-element group 131: 	 branch_block_stmt_31/merge_stmt_108_PhiAck/phi_stmt_109_ack
      -- 
    phi_stmt_109_ack_839_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 131_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_109_ack_0, ack => In_wrap_daemon_CP_0_elements(131)); -- 
    -- CP-element group 132:  transition  bypass 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	84 
    -- CP-element group 132: successors 
    -- CP-element group 132:  members (2) 
      -- CP-element group 132: 	 $exit
      -- CP-element group 132: 	 branch_block_stmt_31/$exit
      -- 
    In_wrap_daemon_CP_0_elements(132) <= In_wrap_daemon_CP_0_elements(84);
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ED_52 : std_logic_vector(0 downto 0);
    signal EQ_u1_u1_117_wire : std_logic_vector(0 downto 0);
    signal EQ_u1_u1_74_wire : std_logic_vector(0 downto 0);
    signal MUX_105_wire : std_logic_vector(14 downto 0);
    signal MUX_99_wire : std_logic_vector(14 downto 0);
    signal RPIPE_w_in_buf_119_wire : std_logic_vector(127 downto 0);
    signal RPIPE_w_in_buf_123_wire : std_logic_vector(127 downto 0);
    signal RPIPE_w_in_buf_148_wire : std_logic_vector(127 downto 0);
    signal R_MAX_COUNT_100_wire_constant : std_logic_vector(14 downto 0);
    signal R_MAX_COUNT_139_wire_constant : std_logic_vector(14 downto 0);
    signal R_MAX_COUNT_157_wire_constant : std_logic_vector(14 downto 0);
    signal R_MAX_COUNT_94_wire_constant : std_logic_vector(14 downto 0);
    signal R_MAX_COUNT_97_wire_constant : std_logic_vector(14 downto 0);
    signal R_ONE_COUNT_111_wire_constant : std_logic_vector(14 downto 0);
    signal UGE_u15_u1_102_wire : std_logic_vector(0 downto 0);
    signal ULT_u15_u1_134_wire : std_logic_vector(0 downto 0);
    signal ULT_u15_u1_140_wire : std_logic_vector(0 downto 0);
    signal ULT_u15_u1_158_wire : std_logic_vector(0 downto 0);
    signal ULT_u15_u1_96_wire : std_logic_vector(0 downto 0);
    signal count_70 : std_logic_vector(14 downto 0);
    signal count_blocks_107 : std_logic_vector(14 downto 0);
    signal count_var2_142 : std_logic_vector(14 downto 0);
    signal count_var_109 : std_logic_vector(14 downto 0);
    signal got_new_key_61 : std_logic_vector(0 downto 0);
    signal head0_38 : std_logic_vector(63 downto 0);
    signal head1_42 : std_logic_vector(63 downto 0);
    signal head_in_34 : std_logic_vector(127 downto 0);
    signal keyA_81 : std_logic_vector(63 downto 0);
    signal keyB_85 : std_logic_vector(63 downto 0);
    signal key_77 : std_logic_vector(127 downto 0);
    signal konst_104_wire_constant : std_logic_vector(14 downto 0);
    signal konst_116_wire_constant : std_logic_vector(0 downto 0);
    signal konst_128_wire_constant : std_logic_vector(14 downto 0);
    signal konst_152_wire_constant : std_logic_vector(14 downto 0);
    signal konst_73_wire_constant : std_logic_vector(0 downto 0);
    signal konst_98_wire_constant : std_logic_vector(14 downto 0);
    signal mode_57 : std_logic_vector(2 downto 0);
    signal n_count_var2_154 : std_logic_vector(14 downto 0);
    signal n_count_var2_154_145_buffered : std_logic_vector(14 downto 0);
    signal n_count_var_130 : std_logic_vector(14 downto 0);
    signal n_count_var_130_112_buffered : std_logic_vector(14 downto 0);
    signal n_count_var_130_144_buffered : std_logic_vector(14 downto 0);
    signal xxIn_wrap_daemonxxMAX_COUNT : std_logic_vector(14 downto 0);
    signal xxIn_wrap_daemonxxONE_COUNT : std_logic_vector(14 downto 0);
    signal xxIn_wrap_daemonxxZERO_COUNT : std_logic_vector(14 downto 0);
    signal xxx_66 : std_logic_vector(43 downto 0);
    -- 
  begin -- 
    R_MAX_COUNT_100_wire_constant <= "000000111111111";
    R_MAX_COUNT_139_wire_constant <= "000000111111111";
    R_MAX_COUNT_157_wire_constant <= "000000111111111";
    R_MAX_COUNT_94_wire_constant <= "000000111111111";
    R_MAX_COUNT_97_wire_constant <= "000000111111111";
    R_ONE_COUNT_111_wire_constant <= "000000000000001";
    konst_104_wire_constant <= "000000000000000";
    konst_116_wire_constant <= "0";
    konst_128_wire_constant <= "000000000000001";
    konst_152_wire_constant <= "000000000000001";
    konst_73_wire_constant <= "1";
    konst_98_wire_constant <= "000000000000000";
    xxIn_wrap_daemonxxMAX_COUNT <= "000000111111111";
    xxIn_wrap_daemonxxONE_COUNT <= "000000000000001";
    xxIn_wrap_daemonxxZERO_COUNT <= "000000000000000";
    phi_stmt_109: Block -- phi operator 
      signal idata: std_logic_vector(29 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ONE_COUNT_111_wire_constant & n_count_var_130_112_buffered;
      req <= phi_stmt_109_req_0 & phi_stmt_109_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_109",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 15) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_109_ack_0,
          idata => idata,
          odata => count_var_109,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_109
    phi_stmt_142: Block -- phi operator 
      signal idata: std_logic_vector(29 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= n_count_var_130_144_buffered & n_count_var2_154_145_buffered;
      req <= phi_stmt_142_req_0 & phi_stmt_142_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_142",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 15) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_142_ack_0,
          idata => idata,
          odata => count_var2_142,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_142
    -- flow-through select operator MUX_105_inst
    MUX_105_wire <= count_70 when (UGE_u15_u1_102_wire(0) /=  '0') else konst_104_wire_constant;
    -- flow-through select operator MUX_99_inst
    MUX_99_wire <= R_MAX_COUNT_97_wire_constant when (ULT_u15_u1_96_wire(0) /=  '0') else konst_98_wire_constant;
    -- flow-through slice operator slice_37_inst
    head0_38 <= head_in_34(127 downto 64);
    -- flow-through slice operator slice_41_inst
    head1_42 <= head_in_34(63 downto 0);
    -- flow-through slice operator slice_51_inst
    ED_52 <= head1_42(63 downto 63);
    -- flow-through slice operator slice_56_inst
    mode_57 <= head1_42(62 downto 60);
    -- flow-through slice operator slice_60_inst
    got_new_key_61 <= head1_42(59 downto 59);
    -- flow-through slice operator slice_65_inst
    xxx_66 <= head1_42(58 downto 15);
    -- flow-through slice operator slice_69_inst
    count_70 <= head1_42(14 downto 0);
    slice_80_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_80_inst_req_0;
      slice_80_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_80_inst_req_1;
      slice_80_inst_ack_1<= update_ack(0);
      slice_80_inst: SliceSplitProtocol generic map(name => "slice_80_inst", in_data_width => 128, high_index => 127, low_index => 64, buffering => 1, flow_through => false,  full_rate => false) -- 
        port map( din => key_77, dout => keyA_81, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_84_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_84_inst_req_0;
      slice_84_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_84_inst_req_1;
      slice_84_inst_ack_1<= update_ack(0);
      slice_84_inst: SliceSplitProtocol generic map(name => "slice_84_inst", in_data_width => 128, high_index => 63, low_index => 0, buffering => 1, flow_through => false,  full_rate => false) -- 
        port map( din => key_77, dout => keyB_85, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    n_count_var2_154_145_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_count_var2_154_145_buf_req_0;
      n_count_var2_154_145_buf_ack_0<= wack(0);
      rreq(0) <= n_count_var2_154_145_buf_req_1;
      n_count_var2_154_145_buf_ack_1<= rack(0);
      n_count_var2_154_145_buf : InterlockBuffer generic map ( -- 
        name => "n_count_var2_154_145_buf",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 15,
        out_data_width => 15,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_count_var2_154,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_count_var2_154_145_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_count_var_130_112_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_count_var_130_112_buf_req_0;
      n_count_var_130_112_buf_ack_0<= wack(0);
      rreq(0) <= n_count_var_130_112_buf_req_1;
      n_count_var_130_112_buf_ack_1<= rack(0);
      n_count_var_130_112_buf : InterlockBuffer generic map ( -- 
        name => "n_count_var_130_112_buf",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 15,
        out_data_width => 15,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_count_var_130,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_count_var_130_112_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_count_var_130_144_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_count_var_130_144_buf_req_0;
      n_count_var_130_144_buf_ack_0<= wack(0);
      rreq(0) <= n_count_var_130_144_buf_req_1;
      n_count_var_130_144_buf_ack_1<= rack(0);
      n_count_var_130_144_buf : InterlockBuffer generic map ( -- 
        name => "n_count_var_130_144_buf",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 15,
        out_data_width => 15,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_count_var_130,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_count_var_130_144_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    if_stmt_114_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= EQ_u1_u1_117_wire;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_114_branch", condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_114_branch_req_0,
          ack0 => if_stmt_114_branch_ack_0,
          ack1 => if_stmt_114_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_131_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= ULT_u15_u1_134_wire;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_131_branch", condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_131_branch_req_0,
          ack0 => if_stmt_131_branch_ack_0,
          ack1 => if_stmt_131_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_137_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= ULT_u15_u1_140_wire;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_137_branch", condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_137_branch_req_0,
          ack0 => if_stmt_137_branch_ack_0,
          ack1 => if_stmt_137_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_155_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= ULT_u15_u1_158_wire;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_155_branch", condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_155_branch_req_0,
          ack0 => if_stmt_155_branch_ack_0,
          ack1 => if_stmt_155_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_71_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= EQ_u1_u1_74_wire;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_71_branch", condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_71_branch_req_0,
          ack0 => if_stmt_71_branch_ack_0,
          ack1 => if_stmt_71_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u15_u15_129_inst
    process(count_var_109) -- 
      variable tmp_var : std_logic_vector(14 downto 0); -- 
    begin -- 
      ApIntAdd_proc(count_var_109, konst_128_wire_constant, tmp_var);
      n_count_var_130 <= tmp_var; -- 
    end process;
    -- binary operator ADD_u15_u15_153_inst
    process(count_var2_142) -- 
      variable tmp_var : std_logic_vector(14 downto 0); -- 
    begin -- 
      ApIntAdd_proc(count_var2_142, konst_152_wire_constant, tmp_var);
      n_count_var2_154 <= tmp_var; -- 
    end process;
    -- binary operator EQ_u1_u1_117_inst
    process(ED_52) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(ED_52, konst_116_wire_constant, tmp_var);
      EQ_u1_u1_117_wire <= tmp_var; -- 
    end process;
    -- binary operator EQ_u1_u1_74_inst
    process(got_new_key_61) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(got_new_key_61, konst_73_wire_constant, tmp_var);
      EQ_u1_u1_74_wire <= tmp_var; -- 
    end process;
    -- shared split operator group (4) : OR_u15_u15_106_inst 
    ApIntOr_group_4: Block -- 
      signal data_in: std_logic_vector(29 downto 0);
      signal data_out: std_logic_vector(14 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= MUX_99_wire & MUX_105_wire;
      count_blocks_107 <= data_out(14 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= OR_u15_u15_106_inst_req_0;
      OR_u15_u15_106_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= OR_u15_u15_106_inst_req_1;
      OR_u15_u15_106_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(name => "gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          name => "ApIntOr_group_4",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 15,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 15, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 15,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 4
    -- binary operator UGE_u15_u1_102_inst
    process(R_MAX_COUNT_100_wire_constant, count_70) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUge_proc(R_MAX_COUNT_100_wire_constant, count_70, tmp_var);
      UGE_u15_u1_102_wire <= tmp_var; -- 
    end process;
    -- binary operator ULT_u15_u1_134_inst
    process(count_var_109, count_blocks_107) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(count_var_109, count_blocks_107, tmp_var);
      ULT_u15_u1_134_wire <= tmp_var; -- 
    end process;
    -- binary operator ULT_u15_u1_140_inst
    process(count_var_109) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(count_var_109, R_MAX_COUNT_139_wire_constant, tmp_var);
      ULT_u15_u1_140_wire <= tmp_var; -- 
    end process;
    -- binary operator ULT_u15_u1_158_inst
    process(count_var2_142) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(count_var2_142, R_MAX_COUNT_157_wire_constant, tmp_var);
      ULT_u15_u1_158_wire <= tmp_var; -- 
    end process;
    -- binary operator ULT_u15_u1_96_inst
    process(R_MAX_COUNT_94_wire_constant, count_70) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(R_MAX_COUNT_94_wire_constant, count_70, tmp_var);
      ULT_u15_u1_96_wire <= tmp_var; -- 
    end process;
    -- shared inport operator group (0) : RPIPE_w_in_buf_148_inst RPIPE_w_in_buf_123_inst RPIPE_w_in_buf_119_inst RPIPE_w_in_buf_33_inst RPIPE_w_in_buf_76_inst 
    InportGroup0: Block -- 
      signal data_out: std_logic_vector(639 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 4 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 4 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 4 downto 0);
      signal guard_vector : std_logic_vector( 4 downto 0);
      constant outBUFs : IntegerArray(4 downto 0) := (4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(4 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false);
      constant guardBuffering: IntegerArray(4 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2);
      -- 
    begin -- 
      reqL_unguarded(4) <= RPIPE_w_in_buf_148_inst_req_0;
      reqL_unguarded(3) <= RPIPE_w_in_buf_123_inst_req_0;
      reqL_unguarded(2) <= RPIPE_w_in_buf_119_inst_req_0;
      reqL_unguarded(1) <= RPIPE_w_in_buf_33_inst_req_0;
      reqL_unguarded(0) <= RPIPE_w_in_buf_76_inst_req_0;
      RPIPE_w_in_buf_148_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_w_in_buf_123_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_w_in_buf_119_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_w_in_buf_33_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_w_in_buf_76_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(4) <= RPIPE_w_in_buf_148_inst_req_1;
      reqR_unguarded(3) <= RPIPE_w_in_buf_123_inst_req_1;
      reqR_unguarded(2) <= RPIPE_w_in_buf_119_inst_req_1;
      reqR_unguarded(1) <= RPIPE_w_in_buf_33_inst_req_1;
      reqR_unguarded(0) <= RPIPE_w_in_buf_76_inst_req_1;
      RPIPE_w_in_buf_148_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_w_in_buf_123_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_w_in_buf_119_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_w_in_buf_33_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_w_in_buf_76_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      gI: SplitGuardInterface generic map(name => "gI", nreqs => 5, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      RPIPE_w_in_buf_148_wire <= data_out(639 downto 512);
      RPIPE_w_in_buf_123_wire <= data_out(511 downto 384);
      RPIPE_w_in_buf_119_wire <= data_out(383 downto 256);
      head_in_34 <= data_out(255 downto 128);
      key_77 <= data_out(127 downto 0);
      w_in_buf_read_0: InputPortRevised -- 
        generic map ( name => "w_in_buf_read_0", data_width => 128,  num_reqs => 5,  output_buffering => outBUFs,   no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => w_in_buf_pipe_read_req(0),
          oack => w_in_buf_pipe_read_ack(0),
          odata => w_in_buf_pipe_read_data(127 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_cmd_in_43_inst WPIPE_cmd_in_86_inst WPIPE_cmd_in_89_inst 
    OutportGroup0: Block -- 
      signal data_in: std_logic_vector(191 downto 0);
      signal sample_req, sample_ack : BooleanArray( 2 downto 0);
      signal update_req, update_ack : BooleanArray( 2 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 2 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 2 downto 0);
      signal guard_vector : std_logic_vector( 2 downto 0);
      constant inBUFs : IntegerArray(2 downto 0) := (2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(2 downto 0) := (0 => false, 1 => false, 2 => false);
      constant guardBuffering: IntegerArray(2 downto 0)  := (0 => 2, 1 => 2, 2 => 2);
      -- 
    begin -- 
      sample_req_unguarded(2) <= WPIPE_cmd_in_43_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_cmd_in_86_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_cmd_in_89_inst_req_0;
      WPIPE_cmd_in_43_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_cmd_in_86_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_cmd_in_89_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(2) <= WPIPE_cmd_in_43_inst_req_1;
      update_req_unguarded(1) <= WPIPE_cmd_in_86_inst_req_1;
      update_req_unguarded(0) <= WPIPE_cmd_in_89_inst_req_1;
      WPIPE_cmd_in_43_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_cmd_in_86_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_cmd_in_89_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      gI: SplitGuardInterface generic map(name => "gI", nreqs => 3, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      data_in <= head1_42 & keyA_81 & keyB_85;
      cmd_in_write_0: OutputPortRevised -- 
        generic map ( name => "cmd_in", data_width => 64, num_reqs => 3, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => cmd_in_pipe_write_req(0),
          oack => cmd_in_pipe_write_ack(0),
          odata => cmd_in_pipe_write_data(63 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_d_in_buf_122_inst 
    OutportGroup1: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_d_in_buf_122_inst_req_0;
      WPIPE_d_in_buf_122_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_d_in_buf_122_inst_req_1;
      WPIPE_d_in_buf_122_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      gI: SplitGuardInterface generic map(name => "gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      data_in <= RPIPE_w_in_buf_123_wire;
      d_in_buf_write_1: OutputPortRevised -- 
        generic map ( name => "d_in_buf", data_width => 128, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => d_in_buf_pipe_write_req(0),
          oack => d_in_buf_pipe_write_ack(0),
          odata => d_in_buf_pipe_write_data(127 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared outport operator group (2) : WPIPE_e_in_buf_118_inst 
    OutportGroup2: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_e_in_buf_118_inst_req_0;
      WPIPE_e_in_buf_118_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_e_in_buf_118_inst_req_1;
      WPIPE_e_in_buf_118_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      gI: SplitGuardInterface generic map(name => "gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      data_in <= RPIPE_w_in_buf_119_wire;
      e_in_buf_write_2: OutputPortRevised -- 
        generic map ( name => "e_in_buf", data_width => 128, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => e_in_buf_pipe_write_req(0),
          oack => e_in_buf_pipe_write_ack(0),
          odata => e_in_buf_pipe_write_data(127 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 2
    -- shared outport operator group (3) : WPIPE_out_wrap_cmd_46_inst 
    OutportGroup3: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_out_wrap_cmd_46_inst_req_0;
      WPIPE_out_wrap_cmd_46_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_out_wrap_cmd_46_inst_req_1;
      WPIPE_out_wrap_cmd_46_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      gI: SplitGuardInterface generic map(name => "gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      data_in <= head1_42;
      out_wrap_cmd_write_3: OutputPortRevised -- 
        generic map ( name => "out_wrap_cmd", data_width => 64, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => out_wrap_cmd_pipe_write_req(0),
          oack => out_wrap_cmd_pipe_write_ack(0),
          odata => out_wrap_cmd_pipe_write_data(63 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 3
    -- shared outport operator group (4) : WPIPE_out_wrap_data_147_inst 
    OutportGroup4: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_out_wrap_data_147_inst_req_0;
      WPIPE_out_wrap_data_147_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_out_wrap_data_147_inst_req_1;
      WPIPE_out_wrap_data_147_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      gI: SplitGuardInterface generic map(name => "gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      data_in <= RPIPE_w_in_buf_148_wire;
      out_wrap_data_write_4: OutputPortRevised -- 
        generic map ( name => "out_wrap_data", data_width => 128, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => out_wrap_data_pipe_write_req(0),
          oack => out_wrap_data_pipe_write_ack(0),
          odata => out_wrap_data_pipe_write_data(127 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 4
    -- 
  end Block; -- data_path
  -- 
end In_wrap_daemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library work;
use work.ahir_system_global_package.all;
entity Inv_Sbox_1_Volatile is -- 
  port ( -- 
    s_in : in  std_logic_vector(7 downto 0);
    s_out : out  std_logic_vector(7 downto 0)-- 
  );
  -- 
end entity Inv_Sbox_1_Volatile;
architecture Inv_Sbox_1_Volatile_arch of Inv_Sbox_1_Volatile is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector(8-1 downto 0);
  signal default_zero_sig: std_logic;
  -- input port buffer signals
  signal s_in_buffer :  std_logic_vector(7 downto 0);
  -- output port buffer signals
  signal s_out_buffer :  std_logic_vector(7 downto 0);
  -- volatile/operator module components. 
  -- 
begin --  
  -- input handling ------------------------------------------------
  s_in_buffer <= s_in;
  -- output handling  -------------------------------------------------------
  s_out <= s_out_buffer;
  -- the control path --------------------------------------------------
  default_zero_sig <= '0';
  -- volatile module, no control path
  -- the data path
  data_path: Block -- 
    signal BITSEL_u8_u1_1002_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1012_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1022_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1032_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1042_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1052_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1062_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1072_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1082_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1092_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1102_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1112_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1122_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1132_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1142_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1152_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1162_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1172_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1182_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1192_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1202_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1212_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1222_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1232_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1242_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1252_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1262_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1272_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1282_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1292_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1302_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1312_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1322_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1332_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1342_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1352_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1362_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1372_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1382_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1392_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1402_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1412_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1422_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1432_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1442_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1452_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1460_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1468_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1476_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1484_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1492_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1500_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1508_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1516_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1524_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1532_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1540_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1548_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1556_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1564_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1572_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1580_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1588_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1596_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1604_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1612_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1620_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1628_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1636_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1644_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1652_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1660_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1668_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1676_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1684_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1692_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1700_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1708_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1716_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1724_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_172_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1732_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1740_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1748_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1756_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1764_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1772_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1780_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1788_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1796_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1804_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1812_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1820_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1828_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_182_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1836_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1844_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1852_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1860_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1868_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1876_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1884_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1892_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1900_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1908_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1916_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1924_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_192_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1932_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1940_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1948_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1956_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1964_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1972_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1980_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1988_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_1996_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2004_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2012_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2020_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2028_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_202_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2036_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2044_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2052_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2060_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2068_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2076_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2084_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2092_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2100_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2108_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2116_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2124_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_212_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2132_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2140_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2148_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2156_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2164_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2172_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2180_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2188_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2196_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2204_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2212_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2220_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2228_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_222_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2236_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2244_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2252_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2260_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2268_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2276_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2284_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2292_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2300_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2308_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2316_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2324_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_232_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2332_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2340_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2348_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2356_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2364_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2372_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2380_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2388_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2396_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2404_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2412_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2420_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2428_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_242_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2436_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2444_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2452_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2460_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_252_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_262_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_272_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_282_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_292_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_302_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_312_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_322_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_332_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_342_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_352_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_362_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_372_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_382_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_392_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_402_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_412_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_422_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_432_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_442_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_452_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_462_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_472_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_482_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_492_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_502_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_512_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_522_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_532_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_542_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_552_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_562_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_572_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_582_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_592_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_602_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_612_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_622_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_632_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_642_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_652_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_662_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_672_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_682_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_692_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_702_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_712_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_722_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_732_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_742_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_752_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_762_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_772_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_782_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_792_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_802_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_812_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_822_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_832_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_842_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_852_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_862_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_872_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_882_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_892_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_902_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_912_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_922_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_932_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_942_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_952_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_962_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_972_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_982_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_992_wire : std_logic_vector(0 downto 0);
    signal IMA0_178 : std_logic_vector(7 downto 0);
    signal IMA100_1178 : std_logic_vector(7 downto 0);
    signal IMA101_1188 : std_logic_vector(7 downto 0);
    signal IMA102_1198 : std_logic_vector(7 downto 0);
    signal IMA103_1208 : std_logic_vector(7 downto 0);
    signal IMA104_1218 : std_logic_vector(7 downto 0);
    signal IMA105_1228 : std_logic_vector(7 downto 0);
    signal IMA106_1238 : std_logic_vector(7 downto 0);
    signal IMA107_1248 : std_logic_vector(7 downto 0);
    signal IMA108_1258 : std_logic_vector(7 downto 0);
    signal IMA109_1268 : std_logic_vector(7 downto 0);
    signal IMA10_278 : std_logic_vector(7 downto 0);
    signal IMA110_1278 : std_logic_vector(7 downto 0);
    signal IMA111_1288 : std_logic_vector(7 downto 0);
    signal IMA112_1298 : std_logic_vector(7 downto 0);
    signal IMA113_1308 : std_logic_vector(7 downto 0);
    signal IMA114_1318 : std_logic_vector(7 downto 0);
    signal IMA115_1328 : std_logic_vector(7 downto 0);
    signal IMA116_1338 : std_logic_vector(7 downto 0);
    signal IMA117_1348 : std_logic_vector(7 downto 0);
    signal IMA118_1358 : std_logic_vector(7 downto 0);
    signal IMA119_1368 : std_logic_vector(7 downto 0);
    signal IMA11_288 : std_logic_vector(7 downto 0);
    signal IMA120_1378 : std_logic_vector(7 downto 0);
    signal IMA121_1388 : std_logic_vector(7 downto 0);
    signal IMA122_1398 : std_logic_vector(7 downto 0);
    signal IMA123_1408 : std_logic_vector(7 downto 0);
    signal IMA124_1418 : std_logic_vector(7 downto 0);
    signal IMA125_1428 : std_logic_vector(7 downto 0);
    signal IMA126_1438 : std_logic_vector(7 downto 0);
    signal IMA127_1448 : std_logic_vector(7 downto 0);
    signal IMA12_298 : std_logic_vector(7 downto 0);
    signal IMA13_308 : std_logic_vector(7 downto 0);
    signal IMA14_318 : std_logic_vector(7 downto 0);
    signal IMA15_328 : std_logic_vector(7 downto 0);
    signal IMA16_338 : std_logic_vector(7 downto 0);
    signal IMA17_348 : std_logic_vector(7 downto 0);
    signal IMA18_358 : std_logic_vector(7 downto 0);
    signal IMA19_368 : std_logic_vector(7 downto 0);
    signal IMA1_188 : std_logic_vector(7 downto 0);
    signal IMA20_378 : std_logic_vector(7 downto 0);
    signal IMA21_388 : std_logic_vector(7 downto 0);
    signal IMA22_398 : std_logic_vector(7 downto 0);
    signal IMA23_408 : std_logic_vector(7 downto 0);
    signal IMA24_418 : std_logic_vector(7 downto 0);
    signal IMA25_428 : std_logic_vector(7 downto 0);
    signal IMA26_438 : std_logic_vector(7 downto 0);
    signal IMA27_448 : std_logic_vector(7 downto 0);
    signal IMA28_458 : std_logic_vector(7 downto 0);
    signal IMA29_468 : std_logic_vector(7 downto 0);
    signal IMA2_198 : std_logic_vector(7 downto 0);
    signal IMA30_478 : std_logic_vector(7 downto 0);
    signal IMA31_488 : std_logic_vector(7 downto 0);
    signal IMA32_498 : std_logic_vector(7 downto 0);
    signal IMA33_508 : std_logic_vector(7 downto 0);
    signal IMA34_518 : std_logic_vector(7 downto 0);
    signal IMA35_528 : std_logic_vector(7 downto 0);
    signal IMA36_538 : std_logic_vector(7 downto 0);
    signal IMA37_548 : std_logic_vector(7 downto 0);
    signal IMA38_558 : std_logic_vector(7 downto 0);
    signal IMA39_568 : std_logic_vector(7 downto 0);
    signal IMA3_208 : std_logic_vector(7 downto 0);
    signal IMA40_578 : std_logic_vector(7 downto 0);
    signal IMA41_588 : std_logic_vector(7 downto 0);
    signal IMA42_598 : std_logic_vector(7 downto 0);
    signal IMA43_608 : std_logic_vector(7 downto 0);
    signal IMA44_618 : std_logic_vector(7 downto 0);
    signal IMA45_628 : std_logic_vector(7 downto 0);
    signal IMA46_638 : std_logic_vector(7 downto 0);
    signal IMA47_648 : std_logic_vector(7 downto 0);
    signal IMA48_658 : std_logic_vector(7 downto 0);
    signal IMA49_668 : std_logic_vector(7 downto 0);
    signal IMA4_218 : std_logic_vector(7 downto 0);
    signal IMA50_678 : std_logic_vector(7 downto 0);
    signal IMA51_688 : std_logic_vector(7 downto 0);
    signal IMA52_698 : std_logic_vector(7 downto 0);
    signal IMA53_708 : std_logic_vector(7 downto 0);
    signal IMA54_718 : std_logic_vector(7 downto 0);
    signal IMA55_728 : std_logic_vector(7 downto 0);
    signal IMA56_738 : std_logic_vector(7 downto 0);
    signal IMA57_748 : std_logic_vector(7 downto 0);
    signal IMA58_758 : std_logic_vector(7 downto 0);
    signal IMA59_768 : std_logic_vector(7 downto 0);
    signal IMA5_228 : std_logic_vector(7 downto 0);
    signal IMA60_778 : std_logic_vector(7 downto 0);
    signal IMA61_788 : std_logic_vector(7 downto 0);
    signal IMA62_798 : std_logic_vector(7 downto 0);
    signal IMA63_808 : std_logic_vector(7 downto 0);
    signal IMA64_818 : std_logic_vector(7 downto 0);
    signal IMA65_828 : std_logic_vector(7 downto 0);
    signal IMA66_838 : std_logic_vector(7 downto 0);
    signal IMA67_848 : std_logic_vector(7 downto 0);
    signal IMA68_858 : std_logic_vector(7 downto 0);
    signal IMA69_868 : std_logic_vector(7 downto 0);
    signal IMA6_238 : std_logic_vector(7 downto 0);
    signal IMA70_878 : std_logic_vector(7 downto 0);
    signal IMA71_888 : std_logic_vector(7 downto 0);
    signal IMA72_898 : std_logic_vector(7 downto 0);
    signal IMA73_908 : std_logic_vector(7 downto 0);
    signal IMA74_918 : std_logic_vector(7 downto 0);
    signal IMA75_928 : std_logic_vector(7 downto 0);
    signal IMA76_938 : std_logic_vector(7 downto 0);
    signal IMA77_948 : std_logic_vector(7 downto 0);
    signal IMA78_958 : std_logic_vector(7 downto 0);
    signal IMA79_968 : std_logic_vector(7 downto 0);
    signal IMA7_248 : std_logic_vector(7 downto 0);
    signal IMA80_978 : std_logic_vector(7 downto 0);
    signal IMA81_988 : std_logic_vector(7 downto 0);
    signal IMA82_998 : std_logic_vector(7 downto 0);
    signal IMA83_1008 : std_logic_vector(7 downto 0);
    signal IMA84_1018 : std_logic_vector(7 downto 0);
    signal IMA85_1028 : std_logic_vector(7 downto 0);
    signal IMA86_1038 : std_logic_vector(7 downto 0);
    signal IMA87_1048 : std_logic_vector(7 downto 0);
    signal IMA88_1058 : std_logic_vector(7 downto 0);
    signal IMA89_1068 : std_logic_vector(7 downto 0);
    signal IMA8_258 : std_logic_vector(7 downto 0);
    signal IMA90_1078 : std_logic_vector(7 downto 0);
    signal IMA91_1088 : std_logic_vector(7 downto 0);
    signal IMA92_1098 : std_logic_vector(7 downto 0);
    signal IMA93_1108 : std_logic_vector(7 downto 0);
    signal IMA94_1118 : std_logic_vector(7 downto 0);
    signal IMA95_1128 : std_logic_vector(7 downto 0);
    signal IMA96_1138 : std_logic_vector(7 downto 0);
    signal IMA97_1148 : std_logic_vector(7 downto 0);
    signal IMA98_1158 : std_logic_vector(7 downto 0);
    signal IMA99_1168 : std_logic_vector(7 downto 0);
    signal IMA9_268 : std_logic_vector(7 downto 0);
    signal IMB0_1456 : std_logic_vector(7 downto 0);
    signal IMB10_1536 : std_logic_vector(7 downto 0);
    signal IMB11_1544 : std_logic_vector(7 downto 0);
    signal IMB12_1552 : std_logic_vector(7 downto 0);
    signal IMB13_1560 : std_logic_vector(7 downto 0);
    signal IMB14_1568 : std_logic_vector(7 downto 0);
    signal IMB15_1576 : std_logic_vector(7 downto 0);
    signal IMB16_1584 : std_logic_vector(7 downto 0);
    signal IMB17_1592 : std_logic_vector(7 downto 0);
    signal IMB18_1600 : std_logic_vector(7 downto 0);
    signal IMB19_1608 : std_logic_vector(7 downto 0);
    signal IMB1_1464 : std_logic_vector(7 downto 0);
    signal IMB20_1616 : std_logic_vector(7 downto 0);
    signal IMB21_1624 : std_logic_vector(7 downto 0);
    signal IMB22_1632 : std_logic_vector(7 downto 0);
    signal IMB23_1640 : std_logic_vector(7 downto 0);
    signal IMB24_1648 : std_logic_vector(7 downto 0);
    signal IMB25_1656 : std_logic_vector(7 downto 0);
    signal IMB26_1664 : std_logic_vector(7 downto 0);
    signal IMB27_1672 : std_logic_vector(7 downto 0);
    signal IMB28_1680 : std_logic_vector(7 downto 0);
    signal IMB29_1688 : std_logic_vector(7 downto 0);
    signal IMB2_1472 : std_logic_vector(7 downto 0);
    signal IMB30_1696 : std_logic_vector(7 downto 0);
    signal IMB31_1704 : std_logic_vector(7 downto 0);
    signal IMB32_1712 : std_logic_vector(7 downto 0);
    signal IMB33_1720 : std_logic_vector(7 downto 0);
    signal IMB34_1728 : std_logic_vector(7 downto 0);
    signal IMB35_1736 : std_logic_vector(7 downto 0);
    signal IMB36_1744 : std_logic_vector(7 downto 0);
    signal IMB37_1752 : std_logic_vector(7 downto 0);
    signal IMB38_1760 : std_logic_vector(7 downto 0);
    signal IMB39_1768 : std_logic_vector(7 downto 0);
    signal IMB3_1480 : std_logic_vector(7 downto 0);
    signal IMB40_1776 : std_logic_vector(7 downto 0);
    signal IMB41_1784 : std_logic_vector(7 downto 0);
    signal IMB42_1792 : std_logic_vector(7 downto 0);
    signal IMB43_1800 : std_logic_vector(7 downto 0);
    signal IMB44_1808 : std_logic_vector(7 downto 0);
    signal IMB45_1816 : std_logic_vector(7 downto 0);
    signal IMB46_1824 : std_logic_vector(7 downto 0);
    signal IMB47_1832 : std_logic_vector(7 downto 0);
    signal IMB48_1840 : std_logic_vector(7 downto 0);
    signal IMB49_1848 : std_logic_vector(7 downto 0);
    signal IMB4_1488 : std_logic_vector(7 downto 0);
    signal IMB50_1856 : std_logic_vector(7 downto 0);
    signal IMB51_1864 : std_logic_vector(7 downto 0);
    signal IMB52_1872 : std_logic_vector(7 downto 0);
    signal IMB53_1880 : std_logic_vector(7 downto 0);
    signal IMB54_1888 : std_logic_vector(7 downto 0);
    signal IMB55_1896 : std_logic_vector(7 downto 0);
    signal IMB56_1904 : std_logic_vector(7 downto 0);
    signal IMB57_1912 : std_logic_vector(7 downto 0);
    signal IMB58_1920 : std_logic_vector(7 downto 0);
    signal IMB59_1928 : std_logic_vector(7 downto 0);
    signal IMB5_1496 : std_logic_vector(7 downto 0);
    signal IMB60_1936 : std_logic_vector(7 downto 0);
    signal IMB61_1944 : std_logic_vector(7 downto 0);
    signal IMB62_1952 : std_logic_vector(7 downto 0);
    signal IMB63_1960 : std_logic_vector(7 downto 0);
    signal IMB6_1504 : std_logic_vector(7 downto 0);
    signal IMB7_1512 : std_logic_vector(7 downto 0);
    signal IMB8_1520 : std_logic_vector(7 downto 0);
    signal IMB9_1528 : std_logic_vector(7 downto 0);
    signal IMC0_1968 : std_logic_vector(7 downto 0);
    signal IMC10_2048 : std_logic_vector(7 downto 0);
    signal IMC11_2056 : std_logic_vector(7 downto 0);
    signal IMC12_2064 : std_logic_vector(7 downto 0);
    signal IMC13_2072 : std_logic_vector(7 downto 0);
    signal IMC14_2080 : std_logic_vector(7 downto 0);
    signal IMC15_2088 : std_logic_vector(7 downto 0);
    signal IMC16_2096 : std_logic_vector(7 downto 0);
    signal IMC17_2104 : std_logic_vector(7 downto 0);
    signal IMC18_2112 : std_logic_vector(7 downto 0);
    signal IMC19_2120 : std_logic_vector(7 downto 0);
    signal IMC1_1976 : std_logic_vector(7 downto 0);
    signal IMC20_2128 : std_logic_vector(7 downto 0);
    signal IMC21_2136 : std_logic_vector(7 downto 0);
    signal IMC22_2144 : std_logic_vector(7 downto 0);
    signal IMC23_2152 : std_logic_vector(7 downto 0);
    signal IMC24_2160 : std_logic_vector(7 downto 0);
    signal IMC25_2168 : std_logic_vector(7 downto 0);
    signal IMC26_2176 : std_logic_vector(7 downto 0);
    signal IMC27_2184 : std_logic_vector(7 downto 0);
    signal IMC28_2192 : std_logic_vector(7 downto 0);
    signal IMC29_2200 : std_logic_vector(7 downto 0);
    signal IMC2_1984 : std_logic_vector(7 downto 0);
    signal IMC30_2208 : std_logic_vector(7 downto 0);
    signal IMC31_2216 : std_logic_vector(7 downto 0);
    signal IMC3_1992 : std_logic_vector(7 downto 0);
    signal IMC4_2000 : std_logic_vector(7 downto 0);
    signal IMC5_2008 : std_logic_vector(7 downto 0);
    signal IMC6_2016 : std_logic_vector(7 downto 0);
    signal IMC7_2024 : std_logic_vector(7 downto 0);
    signal IMC8_2032 : std_logic_vector(7 downto 0);
    signal IMC9_2040 : std_logic_vector(7 downto 0);
    signal IMD0_2224 : std_logic_vector(7 downto 0);
    signal IMD10_2304 : std_logic_vector(7 downto 0);
    signal IMD11_2312 : std_logic_vector(7 downto 0);
    signal IMD12_2320 : std_logic_vector(7 downto 0);
    signal IMD13_2328 : std_logic_vector(7 downto 0);
    signal IMD14_2336 : std_logic_vector(7 downto 0);
    signal IMD15_2344 : std_logic_vector(7 downto 0);
    signal IMD1_2232 : std_logic_vector(7 downto 0);
    signal IMD2_2240 : std_logic_vector(7 downto 0);
    signal IMD3_2248 : std_logic_vector(7 downto 0);
    signal IMD4_2256 : std_logic_vector(7 downto 0);
    signal IMD5_2264 : std_logic_vector(7 downto 0);
    signal IMD6_2272 : std_logic_vector(7 downto 0);
    signal IMD7_2280 : std_logic_vector(7 downto 0);
    signal IMD8_2288 : std_logic_vector(7 downto 0);
    signal IMD9_2296 : std_logic_vector(7 downto 0);
    signal IME0_2352 : std_logic_vector(7 downto 0);
    signal IME1_2360 : std_logic_vector(7 downto 0);
    signal IME2_2368 : std_logic_vector(7 downto 0);
    signal IME3_2376 : std_logic_vector(7 downto 0);
    signal IME4_2384 : std_logic_vector(7 downto 0);
    signal IME5_2392 : std_logic_vector(7 downto 0);
    signal IME6_2400 : std_logic_vector(7 downto 0);
    signal IME7_2408 : std_logic_vector(7 downto 0);
    signal IMF0_2416 : std_logic_vector(7 downto 0);
    signal IMF1_2424 : std_logic_vector(7 downto 0);
    signal IMF2_2432 : std_logic_vector(7 downto 0);
    signal IMF3_2440 : std_logic_vector(7 downto 0);
    signal IMG0_2448 : std_logic_vector(7 downto 0);
    signal IMG1_2456 : std_logic_vector(7 downto 0);
    signal konst_1001_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1011_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1021_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1031_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1041_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1051_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1061_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1071_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1081_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1091_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1101_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1111_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1121_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1131_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1141_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1151_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1161_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1171_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1181_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1191_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1201_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1211_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1221_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1231_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1241_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1251_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1261_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1271_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1281_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1291_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1301_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1311_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1321_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1331_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1341_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1351_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1361_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1371_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1381_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1391_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1401_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1411_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1421_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1431_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1441_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1451_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1459_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1467_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1475_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1483_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1491_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1499_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1507_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1515_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1523_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1531_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1539_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1547_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1555_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1563_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1571_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1579_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1587_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1595_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1603_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1611_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1619_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1627_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1635_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1643_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1651_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1659_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1667_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1675_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1683_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1691_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1699_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1707_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1715_wire_constant : std_logic_vector(7 downto 0);
    signal konst_171_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1723_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1731_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1739_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1747_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1755_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1763_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1771_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1779_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1787_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1795_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1803_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1811_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1819_wire_constant : std_logic_vector(7 downto 0);
    signal konst_181_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1827_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1835_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1843_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1851_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1859_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1867_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1875_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1883_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1891_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1899_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1907_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1915_wire_constant : std_logic_vector(7 downto 0);
    signal konst_191_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1923_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1931_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1939_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1947_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1955_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1963_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1971_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1979_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1987_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1995_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2003_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2011_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2019_wire_constant : std_logic_vector(7 downto 0);
    signal konst_201_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2027_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2035_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2043_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2051_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2059_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2067_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2075_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2083_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2091_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2099_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2107_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2115_wire_constant : std_logic_vector(7 downto 0);
    signal konst_211_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2123_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2131_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2139_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2147_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2155_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2163_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2171_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2179_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2187_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2195_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2203_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2211_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2219_wire_constant : std_logic_vector(7 downto 0);
    signal konst_221_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2227_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2235_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2243_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2251_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2259_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2267_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2275_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2283_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2291_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2299_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2307_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2315_wire_constant : std_logic_vector(7 downto 0);
    signal konst_231_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2323_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2331_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2339_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2347_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2355_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2363_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2371_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2379_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2387_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2395_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2403_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2411_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2419_wire_constant : std_logic_vector(7 downto 0);
    signal konst_241_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2427_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2435_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2443_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2451_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2459_wire_constant : std_logic_vector(7 downto 0);
    signal konst_251_wire_constant : std_logic_vector(7 downto 0);
    signal konst_261_wire_constant : std_logic_vector(7 downto 0);
    signal konst_271_wire_constant : std_logic_vector(7 downto 0);
    signal konst_281_wire_constant : std_logic_vector(7 downto 0);
    signal konst_291_wire_constant : std_logic_vector(7 downto 0);
    signal konst_301_wire_constant : std_logic_vector(7 downto 0);
    signal konst_311_wire_constant : std_logic_vector(7 downto 0);
    signal konst_321_wire_constant : std_logic_vector(7 downto 0);
    signal konst_331_wire_constant : std_logic_vector(7 downto 0);
    signal konst_341_wire_constant : std_logic_vector(7 downto 0);
    signal konst_351_wire_constant : std_logic_vector(7 downto 0);
    signal konst_361_wire_constant : std_logic_vector(7 downto 0);
    signal konst_371_wire_constant : std_logic_vector(7 downto 0);
    signal konst_381_wire_constant : std_logic_vector(7 downto 0);
    signal konst_391_wire_constant : std_logic_vector(7 downto 0);
    signal konst_401_wire_constant : std_logic_vector(7 downto 0);
    signal konst_411_wire_constant : std_logic_vector(7 downto 0);
    signal konst_421_wire_constant : std_logic_vector(7 downto 0);
    signal konst_431_wire_constant : std_logic_vector(7 downto 0);
    signal konst_441_wire_constant : std_logic_vector(7 downto 0);
    signal konst_451_wire_constant : std_logic_vector(7 downto 0);
    signal konst_461_wire_constant : std_logic_vector(7 downto 0);
    signal konst_471_wire_constant : std_logic_vector(7 downto 0);
    signal konst_481_wire_constant : std_logic_vector(7 downto 0);
    signal konst_491_wire_constant : std_logic_vector(7 downto 0);
    signal konst_501_wire_constant : std_logic_vector(7 downto 0);
    signal konst_511_wire_constant : std_logic_vector(7 downto 0);
    signal konst_521_wire_constant : std_logic_vector(7 downto 0);
    signal konst_531_wire_constant : std_logic_vector(7 downto 0);
    signal konst_541_wire_constant : std_logic_vector(7 downto 0);
    signal konst_551_wire_constant : std_logic_vector(7 downto 0);
    signal konst_561_wire_constant : std_logic_vector(7 downto 0);
    signal konst_571_wire_constant : std_logic_vector(7 downto 0);
    signal konst_581_wire_constant : std_logic_vector(7 downto 0);
    signal konst_591_wire_constant : std_logic_vector(7 downto 0);
    signal konst_601_wire_constant : std_logic_vector(7 downto 0);
    signal konst_611_wire_constant : std_logic_vector(7 downto 0);
    signal konst_621_wire_constant : std_logic_vector(7 downto 0);
    signal konst_631_wire_constant : std_logic_vector(7 downto 0);
    signal konst_641_wire_constant : std_logic_vector(7 downto 0);
    signal konst_651_wire_constant : std_logic_vector(7 downto 0);
    signal konst_661_wire_constant : std_logic_vector(7 downto 0);
    signal konst_671_wire_constant : std_logic_vector(7 downto 0);
    signal konst_681_wire_constant : std_logic_vector(7 downto 0);
    signal konst_691_wire_constant : std_logic_vector(7 downto 0);
    signal konst_701_wire_constant : std_logic_vector(7 downto 0);
    signal konst_711_wire_constant : std_logic_vector(7 downto 0);
    signal konst_721_wire_constant : std_logic_vector(7 downto 0);
    signal konst_731_wire_constant : std_logic_vector(7 downto 0);
    signal konst_741_wire_constant : std_logic_vector(7 downto 0);
    signal konst_751_wire_constant : std_logic_vector(7 downto 0);
    signal konst_761_wire_constant : std_logic_vector(7 downto 0);
    signal konst_771_wire_constant : std_logic_vector(7 downto 0);
    signal konst_781_wire_constant : std_logic_vector(7 downto 0);
    signal konst_791_wire_constant : std_logic_vector(7 downto 0);
    signal konst_801_wire_constant : std_logic_vector(7 downto 0);
    signal konst_811_wire_constant : std_logic_vector(7 downto 0);
    signal konst_821_wire_constant : std_logic_vector(7 downto 0);
    signal konst_831_wire_constant : std_logic_vector(7 downto 0);
    signal konst_841_wire_constant : std_logic_vector(7 downto 0);
    signal konst_851_wire_constant : std_logic_vector(7 downto 0);
    signal konst_861_wire_constant : std_logic_vector(7 downto 0);
    signal konst_871_wire_constant : std_logic_vector(7 downto 0);
    signal konst_881_wire_constant : std_logic_vector(7 downto 0);
    signal konst_891_wire_constant : std_logic_vector(7 downto 0);
    signal konst_901_wire_constant : std_logic_vector(7 downto 0);
    signal konst_911_wire_constant : std_logic_vector(7 downto 0);
    signal konst_921_wire_constant : std_logic_vector(7 downto 0);
    signal konst_931_wire_constant : std_logic_vector(7 downto 0);
    signal konst_941_wire_constant : std_logic_vector(7 downto 0);
    signal konst_951_wire_constant : std_logic_vector(7 downto 0);
    signal konst_961_wire_constant : std_logic_vector(7 downto 0);
    signal konst_971_wire_constant : std_logic_vector(7 downto 0);
    signal konst_981_wire_constant : std_logic_vector(7 downto 0);
    signal konst_991_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1004_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1006_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1014_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1016_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1024_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1026_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1034_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1036_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1044_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1046_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1054_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1056_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1064_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1066_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1074_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1076_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1084_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1086_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1094_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1096_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1104_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1106_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1114_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1116_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1124_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1126_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1134_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1136_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1144_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1146_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1154_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1156_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1164_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1166_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1174_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1176_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1184_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1186_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1194_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1196_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1204_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1206_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1214_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1216_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1224_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1226_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1234_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1236_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1244_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1246_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1254_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1256_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1264_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1266_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1274_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1276_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1284_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1286_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1294_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1296_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1304_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1306_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1314_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1316_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1324_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1326_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1334_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1336_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1344_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1346_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1354_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1356_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1364_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1366_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1374_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1376_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1384_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1386_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1394_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1396_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1404_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1406_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1414_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1416_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1424_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1426_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1434_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1436_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1444_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1446_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_174_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_176_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_184_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_186_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_194_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_196_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_204_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_206_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_214_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_216_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_224_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_226_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_234_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_236_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_244_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_246_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_254_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_256_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_264_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_266_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_274_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_276_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_284_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_286_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_294_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_296_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_304_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_306_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_314_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_316_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_324_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_326_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_334_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_336_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_344_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_346_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_354_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_356_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_364_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_366_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_374_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_376_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_384_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_386_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_394_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_396_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_404_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_406_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_414_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_416_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_424_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_426_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_434_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_436_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_444_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_446_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_454_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_456_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_464_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_466_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_474_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_476_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_484_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_486_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_494_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_496_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_504_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_506_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_514_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_516_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_524_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_526_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_534_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_536_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_544_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_546_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_554_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_556_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_564_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_566_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_574_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_576_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_584_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_586_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_594_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_596_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_604_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_606_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_614_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_616_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_624_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_626_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_634_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_636_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_644_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_646_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_654_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_656_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_664_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_666_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_674_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_676_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_684_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_686_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_694_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_696_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_704_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_706_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_714_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_716_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_724_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_726_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_734_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_736_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_744_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_746_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_754_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_756_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_764_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_766_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_774_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_776_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_784_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_786_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_794_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_796_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_804_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_806_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_814_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_816_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_824_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_826_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_834_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_836_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_844_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_846_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_854_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_856_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_864_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_866_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_874_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_876_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_884_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_886_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_894_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_896_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_904_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_906_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_914_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_916_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_924_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_926_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_934_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_936_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_944_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_946_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_954_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_956_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_964_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_966_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_974_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_976_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_984_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_986_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_994_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_996_wire_constant : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    konst_1001_wire_constant <= "00000000";
    konst_1011_wire_constant <= "00000000";
    konst_1021_wire_constant <= "00000000";
    konst_1031_wire_constant <= "00000000";
    konst_1041_wire_constant <= "00000000";
    konst_1051_wire_constant <= "00000000";
    konst_1061_wire_constant <= "00000000";
    konst_1071_wire_constant <= "00000000";
    konst_1081_wire_constant <= "00000000";
    konst_1091_wire_constant <= "00000000";
    konst_1101_wire_constant <= "00000000";
    konst_1111_wire_constant <= "00000000";
    konst_1121_wire_constant <= "00000000";
    konst_1131_wire_constant <= "00000000";
    konst_1141_wire_constant <= "00000000";
    konst_1151_wire_constant <= "00000000";
    konst_1161_wire_constant <= "00000000";
    konst_1171_wire_constant <= "00000000";
    konst_1181_wire_constant <= "00000000";
    konst_1191_wire_constant <= "00000000";
    konst_1201_wire_constant <= "00000000";
    konst_1211_wire_constant <= "00000000";
    konst_1221_wire_constant <= "00000000";
    konst_1231_wire_constant <= "00000000";
    konst_1241_wire_constant <= "00000000";
    konst_1251_wire_constant <= "00000000";
    konst_1261_wire_constant <= "00000000";
    konst_1271_wire_constant <= "00000000";
    konst_1281_wire_constant <= "00000000";
    konst_1291_wire_constant <= "00000000";
    konst_1301_wire_constant <= "00000000";
    konst_1311_wire_constant <= "00000000";
    konst_1321_wire_constant <= "00000000";
    konst_1331_wire_constant <= "00000000";
    konst_1341_wire_constant <= "00000000";
    konst_1351_wire_constant <= "00000000";
    konst_1361_wire_constant <= "00000000";
    konst_1371_wire_constant <= "00000000";
    konst_1381_wire_constant <= "00000000";
    konst_1391_wire_constant <= "00000000";
    konst_1401_wire_constant <= "00000000";
    konst_1411_wire_constant <= "00000000";
    konst_1421_wire_constant <= "00000000";
    konst_1431_wire_constant <= "00000000";
    konst_1441_wire_constant <= "00000000";
    konst_1451_wire_constant <= "00000001";
    konst_1459_wire_constant <= "00000001";
    konst_1467_wire_constant <= "00000001";
    konst_1475_wire_constant <= "00000001";
    konst_1483_wire_constant <= "00000001";
    konst_1491_wire_constant <= "00000001";
    konst_1499_wire_constant <= "00000001";
    konst_1507_wire_constant <= "00000001";
    konst_1515_wire_constant <= "00000001";
    konst_1523_wire_constant <= "00000001";
    konst_1531_wire_constant <= "00000001";
    konst_1539_wire_constant <= "00000001";
    konst_1547_wire_constant <= "00000001";
    konst_1555_wire_constant <= "00000001";
    konst_1563_wire_constant <= "00000001";
    konst_1571_wire_constant <= "00000001";
    konst_1579_wire_constant <= "00000001";
    konst_1587_wire_constant <= "00000001";
    konst_1595_wire_constant <= "00000001";
    konst_1603_wire_constant <= "00000001";
    konst_1611_wire_constant <= "00000001";
    konst_1619_wire_constant <= "00000001";
    konst_1627_wire_constant <= "00000001";
    konst_1635_wire_constant <= "00000001";
    konst_1643_wire_constant <= "00000001";
    konst_1651_wire_constant <= "00000001";
    konst_1659_wire_constant <= "00000001";
    konst_1667_wire_constant <= "00000001";
    konst_1675_wire_constant <= "00000001";
    konst_1683_wire_constant <= "00000001";
    konst_1691_wire_constant <= "00000001";
    konst_1699_wire_constant <= "00000001";
    konst_1707_wire_constant <= "00000001";
    konst_1715_wire_constant <= "00000001";
    konst_171_wire_constant <= "00000000";
    konst_1723_wire_constant <= "00000001";
    konst_1731_wire_constant <= "00000001";
    konst_1739_wire_constant <= "00000001";
    konst_1747_wire_constant <= "00000001";
    konst_1755_wire_constant <= "00000001";
    konst_1763_wire_constant <= "00000001";
    konst_1771_wire_constant <= "00000001";
    konst_1779_wire_constant <= "00000001";
    konst_1787_wire_constant <= "00000001";
    konst_1795_wire_constant <= "00000001";
    konst_1803_wire_constant <= "00000001";
    konst_1811_wire_constant <= "00000001";
    konst_1819_wire_constant <= "00000001";
    konst_181_wire_constant <= "00000000";
    konst_1827_wire_constant <= "00000001";
    konst_1835_wire_constant <= "00000001";
    konst_1843_wire_constant <= "00000001";
    konst_1851_wire_constant <= "00000001";
    konst_1859_wire_constant <= "00000001";
    konst_1867_wire_constant <= "00000001";
    konst_1875_wire_constant <= "00000001";
    konst_1883_wire_constant <= "00000001";
    konst_1891_wire_constant <= "00000001";
    konst_1899_wire_constant <= "00000001";
    konst_1907_wire_constant <= "00000001";
    konst_1915_wire_constant <= "00000001";
    konst_191_wire_constant <= "00000000";
    konst_1923_wire_constant <= "00000001";
    konst_1931_wire_constant <= "00000001";
    konst_1939_wire_constant <= "00000001";
    konst_1947_wire_constant <= "00000001";
    konst_1955_wire_constant <= "00000001";
    konst_1963_wire_constant <= "00000010";
    konst_1971_wire_constant <= "00000010";
    konst_1979_wire_constant <= "00000010";
    konst_1987_wire_constant <= "00000010";
    konst_1995_wire_constant <= "00000010";
    konst_2003_wire_constant <= "00000010";
    konst_2011_wire_constant <= "00000010";
    konst_2019_wire_constant <= "00000010";
    konst_201_wire_constant <= "00000000";
    konst_2027_wire_constant <= "00000010";
    konst_2035_wire_constant <= "00000010";
    konst_2043_wire_constant <= "00000010";
    konst_2051_wire_constant <= "00000010";
    konst_2059_wire_constant <= "00000010";
    konst_2067_wire_constant <= "00000010";
    konst_2075_wire_constant <= "00000010";
    konst_2083_wire_constant <= "00000010";
    konst_2091_wire_constant <= "00000010";
    konst_2099_wire_constant <= "00000010";
    konst_2107_wire_constant <= "00000010";
    konst_2115_wire_constant <= "00000010";
    konst_211_wire_constant <= "00000000";
    konst_2123_wire_constant <= "00000010";
    konst_2131_wire_constant <= "00000010";
    konst_2139_wire_constant <= "00000010";
    konst_2147_wire_constant <= "00000010";
    konst_2155_wire_constant <= "00000010";
    konst_2163_wire_constant <= "00000010";
    konst_2171_wire_constant <= "00000010";
    konst_2179_wire_constant <= "00000010";
    konst_2187_wire_constant <= "00000010";
    konst_2195_wire_constant <= "00000010";
    konst_2203_wire_constant <= "00000010";
    konst_2211_wire_constant <= "00000010";
    konst_2219_wire_constant <= "00000011";
    konst_221_wire_constant <= "00000000";
    konst_2227_wire_constant <= "00000011";
    konst_2235_wire_constant <= "00000011";
    konst_2243_wire_constant <= "00000011";
    konst_2251_wire_constant <= "00000011";
    konst_2259_wire_constant <= "00000011";
    konst_2267_wire_constant <= "00000011";
    konst_2275_wire_constant <= "00000011";
    konst_2283_wire_constant <= "00000011";
    konst_2291_wire_constant <= "00000011";
    konst_2299_wire_constant <= "00000011";
    konst_2307_wire_constant <= "00000011";
    konst_2315_wire_constant <= "00000011";
    konst_231_wire_constant <= "00000000";
    konst_2323_wire_constant <= "00000011";
    konst_2331_wire_constant <= "00000011";
    konst_2339_wire_constant <= "00000011";
    konst_2347_wire_constant <= "00000100";
    konst_2355_wire_constant <= "00000100";
    konst_2363_wire_constant <= "00000100";
    konst_2371_wire_constant <= "00000100";
    konst_2379_wire_constant <= "00000100";
    konst_2387_wire_constant <= "00000100";
    konst_2395_wire_constant <= "00000100";
    konst_2403_wire_constant <= "00000100";
    konst_2411_wire_constant <= "00000101";
    konst_2419_wire_constant <= "00000101";
    konst_241_wire_constant <= "00000000";
    konst_2427_wire_constant <= "00000101";
    konst_2435_wire_constant <= "00000101";
    konst_2443_wire_constant <= "00000110";
    konst_2451_wire_constant <= "00000110";
    konst_2459_wire_constant <= "00000111";
    konst_251_wire_constant <= "00000000";
    konst_261_wire_constant <= "00000000";
    konst_271_wire_constant <= "00000000";
    konst_281_wire_constant <= "00000000";
    konst_291_wire_constant <= "00000000";
    konst_301_wire_constant <= "00000000";
    konst_311_wire_constant <= "00000000";
    konst_321_wire_constant <= "00000000";
    konst_331_wire_constant <= "00000000";
    konst_341_wire_constant <= "00000000";
    konst_351_wire_constant <= "00000000";
    konst_361_wire_constant <= "00000000";
    konst_371_wire_constant <= "00000000";
    konst_381_wire_constant <= "00000000";
    konst_391_wire_constant <= "00000000";
    konst_401_wire_constant <= "00000000";
    konst_411_wire_constant <= "00000000";
    konst_421_wire_constant <= "00000000";
    konst_431_wire_constant <= "00000000";
    konst_441_wire_constant <= "00000000";
    konst_451_wire_constant <= "00000000";
    konst_461_wire_constant <= "00000000";
    konst_471_wire_constant <= "00000000";
    konst_481_wire_constant <= "00000000";
    konst_491_wire_constant <= "00000000";
    konst_501_wire_constant <= "00000000";
    konst_511_wire_constant <= "00000000";
    konst_521_wire_constant <= "00000000";
    konst_531_wire_constant <= "00000000";
    konst_541_wire_constant <= "00000000";
    konst_551_wire_constant <= "00000000";
    konst_561_wire_constant <= "00000000";
    konst_571_wire_constant <= "00000000";
    konst_581_wire_constant <= "00000000";
    konst_591_wire_constant <= "00000000";
    konst_601_wire_constant <= "00000000";
    konst_611_wire_constant <= "00000000";
    konst_621_wire_constant <= "00000000";
    konst_631_wire_constant <= "00000000";
    konst_641_wire_constant <= "00000000";
    konst_651_wire_constant <= "00000000";
    konst_661_wire_constant <= "00000000";
    konst_671_wire_constant <= "00000000";
    konst_681_wire_constant <= "00000000";
    konst_691_wire_constant <= "00000000";
    konst_701_wire_constant <= "00000000";
    konst_711_wire_constant <= "00000000";
    konst_721_wire_constant <= "00000000";
    konst_731_wire_constant <= "00000000";
    konst_741_wire_constant <= "00000000";
    konst_751_wire_constant <= "00000000";
    konst_761_wire_constant <= "00000000";
    konst_771_wire_constant <= "00000000";
    konst_781_wire_constant <= "00000000";
    konst_791_wire_constant <= "00000000";
    konst_801_wire_constant <= "00000000";
    konst_811_wire_constant <= "00000000";
    konst_821_wire_constant <= "00000000";
    konst_831_wire_constant <= "00000000";
    konst_841_wire_constant <= "00000000";
    konst_851_wire_constant <= "00000000";
    konst_861_wire_constant <= "00000000";
    konst_871_wire_constant <= "00000000";
    konst_881_wire_constant <= "00000000";
    konst_891_wire_constant <= "00000000";
    konst_901_wire_constant <= "00000000";
    konst_911_wire_constant <= "00000000";
    konst_921_wire_constant <= "00000000";
    konst_931_wire_constant <= "00000000";
    konst_941_wire_constant <= "00000000";
    konst_951_wire_constant <= "00000000";
    konst_961_wire_constant <= "00000000";
    konst_971_wire_constant <= "00000000";
    konst_981_wire_constant <= "00000000";
    konst_991_wire_constant <= "00000000";
    type_cast_1004_wire_constant <= "10001001";
    type_cast_1006_wire_constant <= "11000101";
    type_cast_1014_wire_constant <= "10110111";
    type_cast_1016_wire_constant <= "01101111";
    type_cast_1024_wire_constant <= "00001110";
    type_cast_1026_wire_constant <= "01100010";
    type_cast_1034_wire_constant <= "00011000";
    type_cast_1036_wire_constant <= "10101010";
    type_cast_1044_wire_constant <= "00011011";
    type_cast_1046_wire_constant <= "10111110";
    type_cast_1054_wire_constant <= "01010110";
    type_cast_1056_wire_constant <= "11111100";
    type_cast_1064_wire_constant <= "01001011";
    type_cast_1066_wire_constant <= "00111110";
    type_cast_1074_wire_constant <= "11010010";
    type_cast_1076_wire_constant <= "11000110";
    type_cast_1084_wire_constant <= "00100000";
    type_cast_1086_wire_constant <= "01111001";
    type_cast_1094_wire_constant <= "11011011";
    type_cast_1096_wire_constant <= "10011010";
    type_cast_1104_wire_constant <= "11111110";
    type_cast_1106_wire_constant <= "11000000";
    type_cast_1114_wire_constant <= "11001101";
    type_cast_1116_wire_constant <= "01111000";
    type_cast_1124_wire_constant <= "11110100";
    type_cast_1126_wire_constant <= "01011010";
    type_cast_1134_wire_constant <= "11011101";
    type_cast_1136_wire_constant <= "00011111";
    type_cast_1144_wire_constant <= "00110011";
    type_cast_1146_wire_constant <= "10101000";
    type_cast_1154_wire_constant <= "00000111";
    type_cast_1156_wire_constant <= "10001000";
    type_cast_1164_wire_constant <= "00110001";
    type_cast_1166_wire_constant <= "11000111";
    type_cast_1174_wire_constant <= "00010010";
    type_cast_1176_wire_constant <= "10110001";
    type_cast_1184_wire_constant <= "01011001";
    type_cast_1186_wire_constant <= "00010000";
    type_cast_1194_wire_constant <= "10000000";
    type_cast_1196_wire_constant <= "00100111";
    type_cast_1204_wire_constant <= "01011111";
    type_cast_1206_wire_constant <= "11101100";
    type_cast_1214_wire_constant <= "01010001";
    type_cast_1216_wire_constant <= "01100000";
    type_cast_1224_wire_constant <= "10101001";
    type_cast_1226_wire_constant <= "01111111";
    type_cast_1234_wire_constant <= "10110101";
    type_cast_1236_wire_constant <= "00011001";
    type_cast_1244_wire_constant <= "00001101";
    type_cast_1246_wire_constant <= "01001010";
    type_cast_1254_wire_constant <= "11100101";
    type_cast_1256_wire_constant <= "00101101";
    type_cast_1264_wire_constant <= "10011111";
    type_cast_1266_wire_constant <= "01111010";
    type_cast_1274_wire_constant <= "11001001";
    type_cast_1276_wire_constant <= "10010011";
    type_cast_1284_wire_constant <= "11101111";
    type_cast_1286_wire_constant <= "10011100";
    type_cast_1294_wire_constant <= "11100000";
    type_cast_1296_wire_constant <= "10100000";
    type_cast_1304_wire_constant <= "01001101";
    type_cast_1306_wire_constant <= "00111011";
    type_cast_1314_wire_constant <= "00101010";
    type_cast_1316_wire_constant <= "10101110";
    type_cast_1324_wire_constant <= "10110000";
    type_cast_1326_wire_constant <= "11110101";
    type_cast_1334_wire_constant <= "11101011";
    type_cast_1336_wire_constant <= "11001000";
    type_cast_1344_wire_constant <= "00111100";
    type_cast_1346_wire_constant <= "10111011";
    type_cast_1354_wire_constant <= "01010011";
    type_cast_1356_wire_constant <= "10000011";
    type_cast_1364_wire_constant <= "01100001";
    type_cast_1366_wire_constant <= "10011001";
    type_cast_1374_wire_constant <= "00101011";
    type_cast_1376_wire_constant <= "00010111";
    type_cast_1384_wire_constant <= "01111110";
    type_cast_1386_wire_constant <= "00000100";
    type_cast_1394_wire_constant <= "01110111";
    type_cast_1396_wire_constant <= "10111010";
    type_cast_1404_wire_constant <= "00100110";
    type_cast_1406_wire_constant <= "11010110";
    type_cast_1414_wire_constant <= "01101001";
    type_cast_1416_wire_constant <= "11100001";
    type_cast_1424_wire_constant <= "01100011";
    type_cast_1426_wire_constant <= "00010100";
    type_cast_1434_wire_constant <= "00100001";
    type_cast_1436_wire_constant <= "01010101";
    type_cast_1444_wire_constant <= "01111101";
    type_cast_1446_wire_constant <= "00001100";
    type_cast_174_wire_constant <= "00001001";
    type_cast_176_wire_constant <= "01010010";
    type_cast_184_wire_constant <= "11010101";
    type_cast_186_wire_constant <= "01101010";
    type_cast_194_wire_constant <= "00110110";
    type_cast_196_wire_constant <= "00110000";
    type_cast_204_wire_constant <= "00111000";
    type_cast_206_wire_constant <= "10100101";
    type_cast_214_wire_constant <= "01000000";
    type_cast_216_wire_constant <= "10111111";
    type_cast_224_wire_constant <= "10011110";
    type_cast_226_wire_constant <= "10100011";
    type_cast_234_wire_constant <= "11110011";
    type_cast_236_wire_constant <= "10000001";
    type_cast_244_wire_constant <= "11111011";
    type_cast_246_wire_constant <= "11010111";
    type_cast_254_wire_constant <= "11100011";
    type_cast_256_wire_constant <= "01111100";
    type_cast_264_wire_constant <= "10000010";
    type_cast_266_wire_constant <= "00111001";
    type_cast_274_wire_constant <= "00101111";
    type_cast_276_wire_constant <= "10011011";
    type_cast_284_wire_constant <= "10000111";
    type_cast_286_wire_constant <= "11111111";
    type_cast_294_wire_constant <= "10001110";
    type_cast_296_wire_constant <= "00110100";
    type_cast_304_wire_constant <= "01000100";
    type_cast_306_wire_constant <= "01000011";
    type_cast_314_wire_constant <= "11011110";
    type_cast_316_wire_constant <= "11000100";
    type_cast_324_wire_constant <= "11001011";
    type_cast_326_wire_constant <= "11101001";
    type_cast_334_wire_constant <= "01111011";
    type_cast_336_wire_constant <= "01010100";
    type_cast_344_wire_constant <= "00110010";
    type_cast_346_wire_constant <= "10010100";
    type_cast_354_wire_constant <= "11000010";
    type_cast_356_wire_constant <= "10100110";
    type_cast_364_wire_constant <= "00111101";
    type_cast_366_wire_constant <= "00100011";
    type_cast_374_wire_constant <= "01001100";
    type_cast_376_wire_constant <= "11101110";
    type_cast_384_wire_constant <= "00001011";
    type_cast_386_wire_constant <= "10010101";
    type_cast_394_wire_constant <= "11111010";
    type_cast_396_wire_constant <= "01000010";
    type_cast_404_wire_constant <= "01001110";
    type_cast_406_wire_constant <= "11000011";
    type_cast_414_wire_constant <= "00101110";
    type_cast_416_wire_constant <= "00001000";
    type_cast_424_wire_constant <= "01100110";
    type_cast_426_wire_constant <= "10100001";
    type_cast_434_wire_constant <= "11011001";
    type_cast_436_wire_constant <= "00101000";
    type_cast_444_wire_constant <= "10110010";
    type_cast_446_wire_constant <= "00100100";
    type_cast_454_wire_constant <= "01011011";
    type_cast_456_wire_constant <= "01110110";
    type_cast_464_wire_constant <= "01001001";
    type_cast_466_wire_constant <= "10100010";
    type_cast_474_wire_constant <= "10001011";
    type_cast_476_wire_constant <= "01101101";
    type_cast_484_wire_constant <= "00100101";
    type_cast_486_wire_constant <= "11010001";
    type_cast_494_wire_constant <= "11111000";
    type_cast_496_wire_constant <= "01110010";
    type_cast_504_wire_constant <= "01100100";
    type_cast_506_wire_constant <= "11110110";
    type_cast_514_wire_constant <= "01101000";
    type_cast_516_wire_constant <= "10000110";
    type_cast_524_wire_constant <= "00010110";
    type_cast_526_wire_constant <= "10011000";
    type_cast_534_wire_constant <= "10100100";
    type_cast_536_wire_constant <= "11010100";
    type_cast_544_wire_constant <= "11001100";
    type_cast_546_wire_constant <= "01011100";
    type_cast_554_wire_constant <= "01100101";
    type_cast_556_wire_constant <= "01011101";
    type_cast_564_wire_constant <= "10010010";
    type_cast_566_wire_constant <= "10110110";
    type_cast_574_wire_constant <= "01110000";
    type_cast_576_wire_constant <= "01101100";
    type_cast_584_wire_constant <= "01010000";
    type_cast_586_wire_constant <= "01001000";
    type_cast_594_wire_constant <= "11101101";
    type_cast_596_wire_constant <= "11111101";
    type_cast_604_wire_constant <= "11011010";
    type_cast_606_wire_constant <= "10111001";
    type_cast_614_wire_constant <= "00010101";
    type_cast_616_wire_constant <= "01011110";
    type_cast_624_wire_constant <= "01010111";
    type_cast_626_wire_constant <= "01000110";
    type_cast_634_wire_constant <= "10001101";
    type_cast_636_wire_constant <= "10100111";
    type_cast_644_wire_constant <= "10000100";
    type_cast_646_wire_constant <= "10011101";
    type_cast_654_wire_constant <= "11011000";
    type_cast_656_wire_constant <= "10010000";
    type_cast_664_wire_constant <= "00000000";
    type_cast_666_wire_constant <= "10101011";
    type_cast_674_wire_constant <= "10111100";
    type_cast_676_wire_constant <= "10001100";
    type_cast_684_wire_constant <= "00001010";
    type_cast_686_wire_constant <= "11010011";
    type_cast_694_wire_constant <= "11100100";
    type_cast_696_wire_constant <= "11110111";
    type_cast_704_wire_constant <= "00000101";
    type_cast_706_wire_constant <= "01011000";
    type_cast_714_wire_constant <= "10110011";
    type_cast_716_wire_constant <= "10111000";
    type_cast_724_wire_constant <= "00000110";
    type_cast_726_wire_constant <= "01000101";
    type_cast_734_wire_constant <= "00101100";
    type_cast_736_wire_constant <= "11010000";
    type_cast_744_wire_constant <= "10001111";
    type_cast_746_wire_constant <= "00011110";
    type_cast_754_wire_constant <= "00111111";
    type_cast_756_wire_constant <= "11001010";
    type_cast_764_wire_constant <= "00000010";
    type_cast_766_wire_constant <= "00001111";
    type_cast_774_wire_constant <= "10101111";
    type_cast_776_wire_constant <= "11000001";
    type_cast_784_wire_constant <= "00000011";
    type_cast_786_wire_constant <= "10111101";
    type_cast_794_wire_constant <= "00010011";
    type_cast_796_wire_constant <= "00000001";
    type_cast_804_wire_constant <= "01101011";
    type_cast_806_wire_constant <= "10001010";
    type_cast_814_wire_constant <= "10010001";
    type_cast_816_wire_constant <= "00111010";
    type_cast_824_wire_constant <= "01000001";
    type_cast_826_wire_constant <= "00010001";
    type_cast_834_wire_constant <= "01100111";
    type_cast_836_wire_constant <= "01001111";
    type_cast_844_wire_constant <= "11101010";
    type_cast_846_wire_constant <= "11011100";
    type_cast_854_wire_constant <= "11110010";
    type_cast_856_wire_constant <= "10010111";
    type_cast_864_wire_constant <= "11001110";
    type_cast_866_wire_constant <= "11001111";
    type_cast_874_wire_constant <= "10110100";
    type_cast_876_wire_constant <= "11110000";
    type_cast_884_wire_constant <= "01110011";
    type_cast_886_wire_constant <= "11100110";
    type_cast_894_wire_constant <= "10101100";
    type_cast_896_wire_constant <= "10010110";
    type_cast_904_wire_constant <= "00100010";
    type_cast_906_wire_constant <= "01110100";
    type_cast_914_wire_constant <= "10101101";
    type_cast_916_wire_constant <= "11100111";
    type_cast_924_wire_constant <= "10000101";
    type_cast_926_wire_constant <= "00110101";
    type_cast_934_wire_constant <= "11111001";
    type_cast_936_wire_constant <= "11100010";
    type_cast_944_wire_constant <= "11101000";
    type_cast_946_wire_constant <= "00110111";
    type_cast_954_wire_constant <= "01110101";
    type_cast_956_wire_constant <= "00011100";
    type_cast_964_wire_constant <= "01101110";
    type_cast_966_wire_constant <= "11011111";
    type_cast_974_wire_constant <= "11110001";
    type_cast_976_wire_constant <= "01000111";
    type_cast_984_wire_constant <= "01110001";
    type_cast_986_wire_constant <= "00011010";
    type_cast_994_wire_constant <= "00101001";
    type_cast_996_wire_constant <= "00011101";
    -- flow-through select operator MUX_1007_inst
    IMA83_1008 <= type_cast_1004_wire_constant when (BITSEL_u8_u1_1002_wire(0) /=  '0') else type_cast_1006_wire_constant;
    -- flow-through select operator MUX_1017_inst
    IMA84_1018 <= type_cast_1014_wire_constant when (BITSEL_u8_u1_1012_wire(0) /=  '0') else type_cast_1016_wire_constant;
    -- flow-through select operator MUX_1027_inst
    IMA85_1028 <= type_cast_1024_wire_constant when (BITSEL_u8_u1_1022_wire(0) /=  '0') else type_cast_1026_wire_constant;
    -- flow-through select operator MUX_1037_inst
    IMA86_1038 <= type_cast_1034_wire_constant when (BITSEL_u8_u1_1032_wire(0) /=  '0') else type_cast_1036_wire_constant;
    -- flow-through select operator MUX_1047_inst
    IMA87_1048 <= type_cast_1044_wire_constant when (BITSEL_u8_u1_1042_wire(0) /=  '0') else type_cast_1046_wire_constant;
    -- flow-through select operator MUX_1057_inst
    IMA88_1058 <= type_cast_1054_wire_constant when (BITSEL_u8_u1_1052_wire(0) /=  '0') else type_cast_1056_wire_constant;
    -- flow-through select operator MUX_1067_inst
    IMA89_1068 <= type_cast_1064_wire_constant when (BITSEL_u8_u1_1062_wire(0) /=  '0') else type_cast_1066_wire_constant;
    -- flow-through select operator MUX_1077_inst
    IMA90_1078 <= type_cast_1074_wire_constant when (BITSEL_u8_u1_1072_wire(0) /=  '0') else type_cast_1076_wire_constant;
    -- flow-through select operator MUX_1087_inst
    IMA91_1088 <= type_cast_1084_wire_constant when (BITSEL_u8_u1_1082_wire(0) /=  '0') else type_cast_1086_wire_constant;
    -- flow-through select operator MUX_1097_inst
    IMA92_1098 <= type_cast_1094_wire_constant when (BITSEL_u8_u1_1092_wire(0) /=  '0') else type_cast_1096_wire_constant;
    -- flow-through select operator MUX_1107_inst
    IMA93_1108 <= type_cast_1104_wire_constant when (BITSEL_u8_u1_1102_wire(0) /=  '0') else type_cast_1106_wire_constant;
    -- flow-through select operator MUX_1117_inst
    IMA94_1118 <= type_cast_1114_wire_constant when (BITSEL_u8_u1_1112_wire(0) /=  '0') else type_cast_1116_wire_constant;
    -- flow-through select operator MUX_1127_inst
    IMA95_1128 <= type_cast_1124_wire_constant when (BITSEL_u8_u1_1122_wire(0) /=  '0') else type_cast_1126_wire_constant;
    -- flow-through select operator MUX_1137_inst
    IMA96_1138 <= type_cast_1134_wire_constant when (BITSEL_u8_u1_1132_wire(0) /=  '0') else type_cast_1136_wire_constant;
    -- flow-through select operator MUX_1147_inst
    IMA97_1148 <= type_cast_1144_wire_constant when (BITSEL_u8_u1_1142_wire(0) /=  '0') else type_cast_1146_wire_constant;
    -- flow-through select operator MUX_1157_inst
    IMA98_1158 <= type_cast_1154_wire_constant when (BITSEL_u8_u1_1152_wire(0) /=  '0') else type_cast_1156_wire_constant;
    -- flow-through select operator MUX_1167_inst
    IMA99_1168 <= type_cast_1164_wire_constant when (BITSEL_u8_u1_1162_wire(0) /=  '0') else type_cast_1166_wire_constant;
    -- flow-through select operator MUX_1177_inst
    IMA100_1178 <= type_cast_1174_wire_constant when (BITSEL_u8_u1_1172_wire(0) /=  '0') else type_cast_1176_wire_constant;
    -- flow-through select operator MUX_1187_inst
    IMA101_1188 <= type_cast_1184_wire_constant when (BITSEL_u8_u1_1182_wire(0) /=  '0') else type_cast_1186_wire_constant;
    -- flow-through select operator MUX_1197_inst
    IMA102_1198 <= type_cast_1194_wire_constant when (BITSEL_u8_u1_1192_wire(0) /=  '0') else type_cast_1196_wire_constant;
    -- flow-through select operator MUX_1207_inst
    IMA103_1208 <= type_cast_1204_wire_constant when (BITSEL_u8_u1_1202_wire(0) /=  '0') else type_cast_1206_wire_constant;
    -- flow-through select operator MUX_1217_inst
    IMA104_1218 <= type_cast_1214_wire_constant when (BITSEL_u8_u1_1212_wire(0) /=  '0') else type_cast_1216_wire_constant;
    -- flow-through select operator MUX_1227_inst
    IMA105_1228 <= type_cast_1224_wire_constant when (BITSEL_u8_u1_1222_wire(0) /=  '0') else type_cast_1226_wire_constant;
    -- flow-through select operator MUX_1237_inst
    IMA106_1238 <= type_cast_1234_wire_constant when (BITSEL_u8_u1_1232_wire(0) /=  '0') else type_cast_1236_wire_constant;
    -- flow-through select operator MUX_1247_inst
    IMA107_1248 <= type_cast_1244_wire_constant when (BITSEL_u8_u1_1242_wire(0) /=  '0') else type_cast_1246_wire_constant;
    -- flow-through select operator MUX_1257_inst
    IMA108_1258 <= type_cast_1254_wire_constant when (BITSEL_u8_u1_1252_wire(0) /=  '0') else type_cast_1256_wire_constant;
    -- flow-through select operator MUX_1267_inst
    IMA109_1268 <= type_cast_1264_wire_constant when (BITSEL_u8_u1_1262_wire(0) /=  '0') else type_cast_1266_wire_constant;
    -- flow-through select operator MUX_1277_inst
    IMA110_1278 <= type_cast_1274_wire_constant when (BITSEL_u8_u1_1272_wire(0) /=  '0') else type_cast_1276_wire_constant;
    -- flow-through select operator MUX_1287_inst
    IMA111_1288 <= type_cast_1284_wire_constant when (BITSEL_u8_u1_1282_wire(0) /=  '0') else type_cast_1286_wire_constant;
    -- flow-through select operator MUX_1297_inst
    IMA112_1298 <= type_cast_1294_wire_constant when (BITSEL_u8_u1_1292_wire(0) /=  '0') else type_cast_1296_wire_constant;
    -- flow-through select operator MUX_1307_inst
    IMA113_1308 <= type_cast_1304_wire_constant when (BITSEL_u8_u1_1302_wire(0) /=  '0') else type_cast_1306_wire_constant;
    -- flow-through select operator MUX_1317_inst
    IMA114_1318 <= type_cast_1314_wire_constant when (BITSEL_u8_u1_1312_wire(0) /=  '0') else type_cast_1316_wire_constant;
    -- flow-through select operator MUX_1327_inst
    IMA115_1328 <= type_cast_1324_wire_constant when (BITSEL_u8_u1_1322_wire(0) /=  '0') else type_cast_1326_wire_constant;
    -- flow-through select operator MUX_1337_inst
    IMA116_1338 <= type_cast_1334_wire_constant when (BITSEL_u8_u1_1332_wire(0) /=  '0') else type_cast_1336_wire_constant;
    -- flow-through select operator MUX_1347_inst
    IMA117_1348 <= type_cast_1344_wire_constant when (BITSEL_u8_u1_1342_wire(0) /=  '0') else type_cast_1346_wire_constant;
    -- flow-through select operator MUX_1357_inst
    IMA118_1358 <= type_cast_1354_wire_constant when (BITSEL_u8_u1_1352_wire(0) /=  '0') else type_cast_1356_wire_constant;
    -- flow-through select operator MUX_1367_inst
    IMA119_1368 <= type_cast_1364_wire_constant when (BITSEL_u8_u1_1362_wire(0) /=  '0') else type_cast_1366_wire_constant;
    -- flow-through select operator MUX_1377_inst
    IMA120_1378 <= type_cast_1374_wire_constant when (BITSEL_u8_u1_1372_wire(0) /=  '0') else type_cast_1376_wire_constant;
    -- flow-through select operator MUX_1387_inst
    IMA121_1388 <= type_cast_1384_wire_constant when (BITSEL_u8_u1_1382_wire(0) /=  '0') else type_cast_1386_wire_constant;
    -- flow-through select operator MUX_1397_inst
    IMA122_1398 <= type_cast_1394_wire_constant when (BITSEL_u8_u1_1392_wire(0) /=  '0') else type_cast_1396_wire_constant;
    -- flow-through select operator MUX_1407_inst
    IMA123_1408 <= type_cast_1404_wire_constant when (BITSEL_u8_u1_1402_wire(0) /=  '0') else type_cast_1406_wire_constant;
    -- flow-through select operator MUX_1417_inst
    IMA124_1418 <= type_cast_1414_wire_constant when (BITSEL_u8_u1_1412_wire(0) /=  '0') else type_cast_1416_wire_constant;
    -- flow-through select operator MUX_1427_inst
    IMA125_1428 <= type_cast_1424_wire_constant when (BITSEL_u8_u1_1422_wire(0) /=  '0') else type_cast_1426_wire_constant;
    -- flow-through select operator MUX_1437_inst
    IMA126_1438 <= type_cast_1434_wire_constant when (BITSEL_u8_u1_1432_wire(0) /=  '0') else type_cast_1436_wire_constant;
    -- flow-through select operator MUX_1447_inst
    IMA127_1448 <= type_cast_1444_wire_constant when (BITSEL_u8_u1_1442_wire(0) /=  '0') else type_cast_1446_wire_constant;
    -- flow-through select operator MUX_1455_inst
    IMB0_1456 <= IMA1_188 when (BITSEL_u8_u1_1452_wire(0) /=  '0') else IMA0_178;
    -- flow-through select operator MUX_1463_inst
    IMB1_1464 <= IMA3_208 when (BITSEL_u8_u1_1460_wire(0) /=  '0') else IMA2_198;
    -- flow-through select operator MUX_1471_inst
    IMB2_1472 <= IMA5_228 when (BITSEL_u8_u1_1468_wire(0) /=  '0') else IMA4_218;
    -- flow-through select operator MUX_1479_inst
    IMB3_1480 <= IMA7_248 when (BITSEL_u8_u1_1476_wire(0) /=  '0') else IMA6_238;
    -- flow-through select operator MUX_1487_inst
    IMB4_1488 <= IMA9_268 when (BITSEL_u8_u1_1484_wire(0) /=  '0') else IMA8_258;
    -- flow-through select operator MUX_1495_inst
    IMB5_1496 <= IMA11_288 when (BITSEL_u8_u1_1492_wire(0) /=  '0') else IMA10_278;
    -- flow-through select operator MUX_1503_inst
    IMB6_1504 <= IMA13_308 when (BITSEL_u8_u1_1500_wire(0) /=  '0') else IMA12_298;
    -- flow-through select operator MUX_1511_inst
    IMB7_1512 <= IMA15_328 when (BITSEL_u8_u1_1508_wire(0) /=  '0') else IMA14_318;
    -- flow-through select operator MUX_1519_inst
    IMB8_1520 <= IMA17_348 when (BITSEL_u8_u1_1516_wire(0) /=  '0') else IMA16_338;
    -- flow-through select operator MUX_1527_inst
    IMB9_1528 <= IMA19_368 when (BITSEL_u8_u1_1524_wire(0) /=  '0') else IMA18_358;
    -- flow-through select operator MUX_1535_inst
    IMB10_1536 <= IMA21_388 when (BITSEL_u8_u1_1532_wire(0) /=  '0') else IMA20_378;
    -- flow-through select operator MUX_1543_inst
    IMB11_1544 <= IMA23_408 when (BITSEL_u8_u1_1540_wire(0) /=  '0') else IMA22_398;
    -- flow-through select operator MUX_1551_inst
    IMB12_1552 <= IMA25_428 when (BITSEL_u8_u1_1548_wire(0) /=  '0') else IMA24_418;
    -- flow-through select operator MUX_1559_inst
    IMB13_1560 <= IMA27_448 when (BITSEL_u8_u1_1556_wire(0) /=  '0') else IMA26_438;
    -- flow-through select operator MUX_1567_inst
    IMB14_1568 <= IMA29_468 when (BITSEL_u8_u1_1564_wire(0) /=  '0') else IMA28_458;
    -- flow-through select operator MUX_1575_inst
    IMB15_1576 <= IMA31_488 when (BITSEL_u8_u1_1572_wire(0) /=  '0') else IMA30_478;
    -- flow-through select operator MUX_1583_inst
    IMB16_1584 <= IMA33_508 when (BITSEL_u8_u1_1580_wire(0) /=  '0') else IMA32_498;
    -- flow-through select operator MUX_1591_inst
    IMB17_1592 <= IMA35_528 when (BITSEL_u8_u1_1588_wire(0) /=  '0') else IMA34_518;
    -- flow-through select operator MUX_1599_inst
    IMB18_1600 <= IMA37_548 when (BITSEL_u8_u1_1596_wire(0) /=  '0') else IMA36_538;
    -- flow-through select operator MUX_1607_inst
    IMB19_1608 <= IMA39_568 when (BITSEL_u8_u1_1604_wire(0) /=  '0') else IMA38_558;
    -- flow-through select operator MUX_1615_inst
    IMB20_1616 <= IMA41_588 when (BITSEL_u8_u1_1612_wire(0) /=  '0') else IMA40_578;
    -- flow-through select operator MUX_1623_inst
    IMB21_1624 <= IMA43_608 when (BITSEL_u8_u1_1620_wire(0) /=  '0') else IMA42_598;
    -- flow-through select operator MUX_1631_inst
    IMB22_1632 <= IMA45_628 when (BITSEL_u8_u1_1628_wire(0) /=  '0') else IMA44_618;
    -- flow-through select operator MUX_1639_inst
    IMB23_1640 <= IMA47_648 when (BITSEL_u8_u1_1636_wire(0) /=  '0') else IMA46_638;
    -- flow-through select operator MUX_1647_inst
    IMB24_1648 <= IMA49_668 when (BITSEL_u8_u1_1644_wire(0) /=  '0') else IMA48_658;
    -- flow-through select operator MUX_1655_inst
    IMB25_1656 <= IMA51_688 when (BITSEL_u8_u1_1652_wire(0) /=  '0') else IMA50_678;
    -- flow-through select operator MUX_1663_inst
    IMB26_1664 <= IMA53_708 when (BITSEL_u8_u1_1660_wire(0) /=  '0') else IMA52_698;
    -- flow-through select operator MUX_1671_inst
    IMB27_1672 <= IMA55_728 when (BITSEL_u8_u1_1668_wire(0) /=  '0') else IMA54_718;
    -- flow-through select operator MUX_1679_inst
    IMB28_1680 <= IMA57_748 when (BITSEL_u8_u1_1676_wire(0) /=  '0') else IMA56_738;
    -- flow-through select operator MUX_1687_inst
    IMB29_1688 <= IMA59_768 when (BITSEL_u8_u1_1684_wire(0) /=  '0') else IMA58_758;
    -- flow-through select operator MUX_1695_inst
    IMB30_1696 <= IMA61_788 when (BITSEL_u8_u1_1692_wire(0) /=  '0') else IMA60_778;
    -- flow-through select operator MUX_1703_inst
    IMB31_1704 <= IMA63_808 when (BITSEL_u8_u1_1700_wire(0) /=  '0') else IMA62_798;
    -- flow-through select operator MUX_1711_inst
    IMB32_1712 <= IMA65_828 when (BITSEL_u8_u1_1708_wire(0) /=  '0') else IMA64_818;
    -- flow-through select operator MUX_1719_inst
    IMB33_1720 <= IMA67_848 when (BITSEL_u8_u1_1716_wire(0) /=  '0') else IMA66_838;
    -- flow-through select operator MUX_1727_inst
    IMB34_1728 <= IMA69_868 when (BITSEL_u8_u1_1724_wire(0) /=  '0') else IMA68_858;
    -- flow-through select operator MUX_1735_inst
    IMB35_1736 <= IMA71_888 when (BITSEL_u8_u1_1732_wire(0) /=  '0') else IMA70_878;
    -- flow-through select operator MUX_1743_inst
    IMB36_1744 <= IMA73_908 when (BITSEL_u8_u1_1740_wire(0) /=  '0') else IMA72_898;
    -- flow-through select operator MUX_1751_inst
    IMB37_1752 <= IMA75_928 when (BITSEL_u8_u1_1748_wire(0) /=  '0') else IMA74_918;
    -- flow-through select operator MUX_1759_inst
    IMB38_1760 <= IMA77_948 when (BITSEL_u8_u1_1756_wire(0) /=  '0') else IMA76_938;
    -- flow-through select operator MUX_1767_inst
    IMB39_1768 <= IMA79_968 when (BITSEL_u8_u1_1764_wire(0) /=  '0') else IMA78_958;
    -- flow-through select operator MUX_1775_inst
    IMB40_1776 <= IMA81_988 when (BITSEL_u8_u1_1772_wire(0) /=  '0') else IMA80_978;
    -- flow-through select operator MUX_177_inst
    IMA0_178 <= type_cast_174_wire_constant when (BITSEL_u8_u1_172_wire(0) /=  '0') else type_cast_176_wire_constant;
    -- flow-through select operator MUX_1783_inst
    IMB41_1784 <= IMA83_1008 when (BITSEL_u8_u1_1780_wire(0) /=  '0') else IMA82_998;
    -- flow-through select operator MUX_1791_inst
    IMB42_1792 <= IMA85_1028 when (BITSEL_u8_u1_1788_wire(0) /=  '0') else IMA84_1018;
    -- flow-through select operator MUX_1799_inst
    IMB43_1800 <= IMA87_1048 when (BITSEL_u8_u1_1796_wire(0) /=  '0') else IMA86_1038;
    -- flow-through select operator MUX_1807_inst
    IMB44_1808 <= IMA89_1068 when (BITSEL_u8_u1_1804_wire(0) /=  '0') else IMA88_1058;
    -- flow-through select operator MUX_1815_inst
    IMB45_1816 <= IMA91_1088 when (BITSEL_u8_u1_1812_wire(0) /=  '0') else IMA90_1078;
    -- flow-through select operator MUX_1823_inst
    IMB46_1824 <= IMA93_1108 when (BITSEL_u8_u1_1820_wire(0) /=  '0') else IMA92_1098;
    -- flow-through select operator MUX_1831_inst
    IMB47_1832 <= IMA95_1128 when (BITSEL_u8_u1_1828_wire(0) /=  '0') else IMA94_1118;
    -- flow-through select operator MUX_1839_inst
    IMB48_1840 <= IMA97_1148 when (BITSEL_u8_u1_1836_wire(0) /=  '0') else IMA96_1138;
    -- flow-through select operator MUX_1847_inst
    IMB49_1848 <= IMA99_1168 when (BITSEL_u8_u1_1844_wire(0) /=  '0') else IMA98_1158;
    -- flow-through select operator MUX_1855_inst
    IMB50_1856 <= IMA101_1188 when (BITSEL_u8_u1_1852_wire(0) /=  '0') else IMA100_1178;
    -- flow-through select operator MUX_1863_inst
    IMB51_1864 <= IMA103_1208 when (BITSEL_u8_u1_1860_wire(0) /=  '0') else IMA102_1198;
    -- flow-through select operator MUX_1871_inst
    IMB52_1872 <= IMA105_1228 when (BITSEL_u8_u1_1868_wire(0) /=  '0') else IMA104_1218;
    -- flow-through select operator MUX_1879_inst
    IMB53_1880 <= IMA107_1248 when (BITSEL_u8_u1_1876_wire(0) /=  '0') else IMA106_1238;
    -- flow-through select operator MUX_187_inst
    IMA1_188 <= type_cast_184_wire_constant when (BITSEL_u8_u1_182_wire(0) /=  '0') else type_cast_186_wire_constant;
    -- flow-through select operator MUX_1887_inst
    IMB54_1888 <= IMA109_1268 when (BITSEL_u8_u1_1884_wire(0) /=  '0') else IMA108_1258;
    -- flow-through select operator MUX_1895_inst
    IMB55_1896 <= IMA111_1288 when (BITSEL_u8_u1_1892_wire(0) /=  '0') else IMA110_1278;
    -- flow-through select operator MUX_1903_inst
    IMB56_1904 <= IMA113_1308 when (BITSEL_u8_u1_1900_wire(0) /=  '0') else IMA112_1298;
    -- flow-through select operator MUX_1911_inst
    IMB57_1912 <= IMA115_1328 when (BITSEL_u8_u1_1908_wire(0) /=  '0') else IMA114_1318;
    -- flow-through select operator MUX_1919_inst
    IMB58_1920 <= IMA117_1348 when (BITSEL_u8_u1_1916_wire(0) /=  '0') else IMA116_1338;
    -- flow-through select operator MUX_1927_inst
    IMB59_1928 <= IMA119_1368 when (BITSEL_u8_u1_1924_wire(0) /=  '0') else IMA118_1358;
    -- flow-through select operator MUX_1935_inst
    IMB60_1936 <= IMA121_1388 when (BITSEL_u8_u1_1932_wire(0) /=  '0') else IMA120_1378;
    -- flow-through select operator MUX_1943_inst
    IMB61_1944 <= IMA123_1408 when (BITSEL_u8_u1_1940_wire(0) /=  '0') else IMA122_1398;
    -- flow-through select operator MUX_1951_inst
    IMB62_1952 <= IMA125_1428 when (BITSEL_u8_u1_1948_wire(0) /=  '0') else IMA124_1418;
    -- flow-through select operator MUX_1959_inst
    IMB63_1960 <= IMA127_1448 when (BITSEL_u8_u1_1956_wire(0) /=  '0') else IMA126_1438;
    -- flow-through select operator MUX_1967_inst
    IMC0_1968 <= IMB1_1464 when (BITSEL_u8_u1_1964_wire(0) /=  '0') else IMB0_1456;
    -- flow-through select operator MUX_1975_inst
    IMC1_1976 <= IMB3_1480 when (BITSEL_u8_u1_1972_wire(0) /=  '0') else IMB2_1472;
    -- flow-through select operator MUX_197_inst
    IMA2_198 <= type_cast_194_wire_constant when (BITSEL_u8_u1_192_wire(0) /=  '0') else type_cast_196_wire_constant;
    -- flow-through select operator MUX_1983_inst
    IMC2_1984 <= IMB5_1496 when (BITSEL_u8_u1_1980_wire(0) /=  '0') else IMB4_1488;
    -- flow-through select operator MUX_1991_inst
    IMC3_1992 <= IMB7_1512 when (BITSEL_u8_u1_1988_wire(0) /=  '0') else IMB6_1504;
    -- flow-through select operator MUX_1999_inst
    IMC4_2000 <= IMB9_1528 when (BITSEL_u8_u1_1996_wire(0) /=  '0') else IMB8_1520;
    -- flow-through select operator MUX_2007_inst
    IMC5_2008 <= IMB11_1544 when (BITSEL_u8_u1_2004_wire(0) /=  '0') else IMB10_1536;
    -- flow-through select operator MUX_2015_inst
    IMC6_2016 <= IMB13_1560 when (BITSEL_u8_u1_2012_wire(0) /=  '0') else IMB12_1552;
    -- flow-through select operator MUX_2023_inst
    IMC7_2024 <= IMB15_1576 when (BITSEL_u8_u1_2020_wire(0) /=  '0') else IMB14_1568;
    -- flow-through select operator MUX_2031_inst
    IMC8_2032 <= IMB17_1592 when (BITSEL_u8_u1_2028_wire(0) /=  '0') else IMB16_1584;
    -- flow-through select operator MUX_2039_inst
    IMC9_2040 <= IMB19_1608 when (BITSEL_u8_u1_2036_wire(0) /=  '0') else IMB18_1600;
    -- flow-through select operator MUX_2047_inst
    IMC10_2048 <= IMB21_1624 when (BITSEL_u8_u1_2044_wire(0) /=  '0') else IMB20_1616;
    -- flow-through select operator MUX_2055_inst
    IMC11_2056 <= IMB23_1640 when (BITSEL_u8_u1_2052_wire(0) /=  '0') else IMB22_1632;
    -- flow-through select operator MUX_2063_inst
    IMC12_2064 <= IMB25_1656 when (BITSEL_u8_u1_2060_wire(0) /=  '0') else IMB24_1648;
    -- flow-through select operator MUX_2071_inst
    IMC13_2072 <= IMB27_1672 when (BITSEL_u8_u1_2068_wire(0) /=  '0') else IMB26_1664;
    -- flow-through select operator MUX_2079_inst
    IMC14_2080 <= IMB29_1688 when (BITSEL_u8_u1_2076_wire(0) /=  '0') else IMB28_1680;
    -- flow-through select operator MUX_207_inst
    IMA3_208 <= type_cast_204_wire_constant when (BITSEL_u8_u1_202_wire(0) /=  '0') else type_cast_206_wire_constant;
    -- flow-through select operator MUX_2087_inst
    IMC15_2088 <= IMB31_1704 when (BITSEL_u8_u1_2084_wire(0) /=  '0') else IMB30_1696;
    -- flow-through select operator MUX_2095_inst
    IMC16_2096 <= IMB33_1720 when (BITSEL_u8_u1_2092_wire(0) /=  '0') else IMB32_1712;
    -- flow-through select operator MUX_2103_inst
    IMC17_2104 <= IMB35_1736 when (BITSEL_u8_u1_2100_wire(0) /=  '0') else IMB34_1728;
    -- flow-through select operator MUX_2111_inst
    IMC18_2112 <= IMB37_1752 when (BITSEL_u8_u1_2108_wire(0) /=  '0') else IMB36_1744;
    -- flow-through select operator MUX_2119_inst
    IMC19_2120 <= IMB39_1768 when (BITSEL_u8_u1_2116_wire(0) /=  '0') else IMB38_1760;
    -- flow-through select operator MUX_2127_inst
    IMC20_2128 <= IMB41_1784 when (BITSEL_u8_u1_2124_wire(0) /=  '0') else IMB40_1776;
    -- flow-through select operator MUX_2135_inst
    IMC21_2136 <= IMB43_1800 when (BITSEL_u8_u1_2132_wire(0) /=  '0') else IMB42_1792;
    -- flow-through select operator MUX_2143_inst
    IMC22_2144 <= IMB45_1816 when (BITSEL_u8_u1_2140_wire(0) /=  '0') else IMB44_1808;
    -- flow-through select operator MUX_2151_inst
    IMC23_2152 <= IMB47_1832 when (BITSEL_u8_u1_2148_wire(0) /=  '0') else IMB46_1824;
    -- flow-through select operator MUX_2159_inst
    IMC24_2160 <= IMB49_1848 when (BITSEL_u8_u1_2156_wire(0) /=  '0') else IMB48_1840;
    -- flow-through select operator MUX_2167_inst
    IMC25_2168 <= IMB51_1864 when (BITSEL_u8_u1_2164_wire(0) /=  '0') else IMB50_1856;
    -- flow-through select operator MUX_2175_inst
    IMC26_2176 <= IMB53_1880 when (BITSEL_u8_u1_2172_wire(0) /=  '0') else IMB52_1872;
    -- flow-through select operator MUX_217_inst
    IMA4_218 <= type_cast_214_wire_constant when (BITSEL_u8_u1_212_wire(0) /=  '0') else type_cast_216_wire_constant;
    -- flow-through select operator MUX_2183_inst
    IMC27_2184 <= IMB55_1896 when (BITSEL_u8_u1_2180_wire(0) /=  '0') else IMB54_1888;
    -- flow-through select operator MUX_2191_inst
    IMC28_2192 <= IMB57_1912 when (BITSEL_u8_u1_2188_wire(0) /=  '0') else IMB56_1904;
    -- flow-through select operator MUX_2199_inst
    IMC29_2200 <= IMB59_1928 when (BITSEL_u8_u1_2196_wire(0) /=  '0') else IMB58_1920;
    -- flow-through select operator MUX_2207_inst
    IMC30_2208 <= IMB61_1944 when (BITSEL_u8_u1_2204_wire(0) /=  '0') else IMB60_1936;
    -- flow-through select operator MUX_2215_inst
    IMC31_2216 <= IMB63_1960 when (BITSEL_u8_u1_2212_wire(0) /=  '0') else IMB62_1952;
    -- flow-through select operator MUX_2223_inst
    IMD0_2224 <= IMC1_1976 when (BITSEL_u8_u1_2220_wire(0) /=  '0') else IMC0_1968;
    -- flow-through select operator MUX_2231_inst
    IMD1_2232 <= IMC3_1992 when (BITSEL_u8_u1_2228_wire(0) /=  '0') else IMC2_1984;
    -- flow-through select operator MUX_2239_inst
    IMD2_2240 <= IMC5_2008 when (BITSEL_u8_u1_2236_wire(0) /=  '0') else IMC4_2000;
    -- flow-through select operator MUX_2247_inst
    IMD3_2248 <= IMC7_2024 when (BITSEL_u8_u1_2244_wire(0) /=  '0') else IMC6_2016;
    -- flow-through select operator MUX_2255_inst
    IMD4_2256 <= IMC9_2040 when (BITSEL_u8_u1_2252_wire(0) /=  '0') else IMC8_2032;
    -- flow-through select operator MUX_2263_inst
    IMD5_2264 <= IMC11_2056 when (BITSEL_u8_u1_2260_wire(0) /=  '0') else IMC10_2048;
    -- flow-through select operator MUX_2271_inst
    IMD6_2272 <= IMC13_2072 when (BITSEL_u8_u1_2268_wire(0) /=  '0') else IMC12_2064;
    -- flow-through select operator MUX_2279_inst
    IMD7_2280 <= IMC15_2088 when (BITSEL_u8_u1_2276_wire(0) /=  '0') else IMC14_2080;
    -- flow-through select operator MUX_227_inst
    IMA5_228 <= type_cast_224_wire_constant when (BITSEL_u8_u1_222_wire(0) /=  '0') else type_cast_226_wire_constant;
    -- flow-through select operator MUX_2287_inst
    IMD8_2288 <= IMC17_2104 when (BITSEL_u8_u1_2284_wire(0) /=  '0') else IMC16_2096;
    -- flow-through select operator MUX_2295_inst
    IMD9_2296 <= IMC19_2120 when (BITSEL_u8_u1_2292_wire(0) /=  '0') else IMC18_2112;
    -- flow-through select operator MUX_2303_inst
    IMD10_2304 <= IMC21_2136 when (BITSEL_u8_u1_2300_wire(0) /=  '0') else IMC20_2128;
    -- flow-through select operator MUX_2311_inst
    IMD11_2312 <= IMC23_2152 when (BITSEL_u8_u1_2308_wire(0) /=  '0') else IMC22_2144;
    -- flow-through select operator MUX_2319_inst
    IMD12_2320 <= IMC25_2168 when (BITSEL_u8_u1_2316_wire(0) /=  '0') else IMC24_2160;
    -- flow-through select operator MUX_2327_inst
    IMD13_2328 <= IMC27_2184 when (BITSEL_u8_u1_2324_wire(0) /=  '0') else IMC26_2176;
    -- flow-through select operator MUX_2335_inst
    IMD14_2336 <= IMC29_2200 when (BITSEL_u8_u1_2332_wire(0) /=  '0') else IMC28_2192;
    -- flow-through select operator MUX_2343_inst
    IMD15_2344 <= IMC31_2216 when (BITSEL_u8_u1_2340_wire(0) /=  '0') else IMC30_2208;
    -- flow-through select operator MUX_2351_inst
    IME0_2352 <= IMD1_2232 when (BITSEL_u8_u1_2348_wire(0) /=  '0') else IMD0_2224;
    -- flow-through select operator MUX_2359_inst
    IME1_2360 <= IMD3_2248 when (BITSEL_u8_u1_2356_wire(0) /=  '0') else IMD2_2240;
    -- flow-through select operator MUX_2367_inst
    IME2_2368 <= IMD5_2264 when (BITSEL_u8_u1_2364_wire(0) /=  '0') else IMD4_2256;
    -- flow-through select operator MUX_2375_inst
    IME3_2376 <= IMD7_2280 when (BITSEL_u8_u1_2372_wire(0) /=  '0') else IMD6_2272;
    -- flow-through select operator MUX_237_inst
    IMA6_238 <= type_cast_234_wire_constant when (BITSEL_u8_u1_232_wire(0) /=  '0') else type_cast_236_wire_constant;
    -- flow-through select operator MUX_2383_inst
    IME4_2384 <= IMD9_2296 when (BITSEL_u8_u1_2380_wire(0) /=  '0') else IMD8_2288;
    -- flow-through select operator MUX_2391_inst
    IME5_2392 <= IMD11_2312 when (BITSEL_u8_u1_2388_wire(0) /=  '0') else IMD10_2304;
    -- flow-through select operator MUX_2399_inst
    IME6_2400 <= IMD13_2328 when (BITSEL_u8_u1_2396_wire(0) /=  '0') else IMD12_2320;
    -- flow-through select operator MUX_2407_inst
    IME7_2408 <= IMD15_2344 when (BITSEL_u8_u1_2404_wire(0) /=  '0') else IMD14_2336;
    -- flow-through select operator MUX_2415_inst
    IMF0_2416 <= IME1_2360 when (BITSEL_u8_u1_2412_wire(0) /=  '0') else IME0_2352;
    -- flow-through select operator MUX_2423_inst
    IMF1_2424 <= IME3_2376 when (BITSEL_u8_u1_2420_wire(0) /=  '0') else IME2_2368;
    -- flow-through select operator MUX_2431_inst
    IMF2_2432 <= IME5_2392 when (BITSEL_u8_u1_2428_wire(0) /=  '0') else IME4_2384;
    -- flow-through select operator MUX_2439_inst
    IMF3_2440 <= IME7_2408 when (BITSEL_u8_u1_2436_wire(0) /=  '0') else IME6_2400;
    -- flow-through select operator MUX_2447_inst
    IMG0_2448 <= IMF1_2424 when (BITSEL_u8_u1_2444_wire(0) /=  '0') else IMF0_2416;
    -- flow-through select operator MUX_2455_inst
    IMG1_2456 <= IMF3_2440 when (BITSEL_u8_u1_2452_wire(0) /=  '0') else IMF2_2432;
    -- flow-through select operator MUX_2463_inst
    s_out_buffer <= IMG1_2456 when (BITSEL_u8_u1_2460_wire(0) /=  '0') else IMG0_2448;
    -- flow-through select operator MUX_247_inst
    IMA7_248 <= type_cast_244_wire_constant when (BITSEL_u8_u1_242_wire(0) /=  '0') else type_cast_246_wire_constant;
    -- flow-through select operator MUX_257_inst
    IMA8_258 <= type_cast_254_wire_constant when (BITSEL_u8_u1_252_wire(0) /=  '0') else type_cast_256_wire_constant;
    -- flow-through select operator MUX_267_inst
    IMA9_268 <= type_cast_264_wire_constant when (BITSEL_u8_u1_262_wire(0) /=  '0') else type_cast_266_wire_constant;
    -- flow-through select operator MUX_277_inst
    IMA10_278 <= type_cast_274_wire_constant when (BITSEL_u8_u1_272_wire(0) /=  '0') else type_cast_276_wire_constant;
    -- flow-through select operator MUX_287_inst
    IMA11_288 <= type_cast_284_wire_constant when (BITSEL_u8_u1_282_wire(0) /=  '0') else type_cast_286_wire_constant;
    -- flow-through select operator MUX_297_inst
    IMA12_298 <= type_cast_294_wire_constant when (BITSEL_u8_u1_292_wire(0) /=  '0') else type_cast_296_wire_constant;
    -- flow-through select operator MUX_307_inst
    IMA13_308 <= type_cast_304_wire_constant when (BITSEL_u8_u1_302_wire(0) /=  '0') else type_cast_306_wire_constant;
    -- flow-through select operator MUX_317_inst
    IMA14_318 <= type_cast_314_wire_constant when (BITSEL_u8_u1_312_wire(0) /=  '0') else type_cast_316_wire_constant;
    -- flow-through select operator MUX_327_inst
    IMA15_328 <= type_cast_324_wire_constant when (BITSEL_u8_u1_322_wire(0) /=  '0') else type_cast_326_wire_constant;
    -- flow-through select operator MUX_337_inst
    IMA16_338 <= type_cast_334_wire_constant when (BITSEL_u8_u1_332_wire(0) /=  '0') else type_cast_336_wire_constant;
    -- flow-through select operator MUX_347_inst
    IMA17_348 <= type_cast_344_wire_constant when (BITSEL_u8_u1_342_wire(0) /=  '0') else type_cast_346_wire_constant;
    -- flow-through select operator MUX_357_inst
    IMA18_358 <= type_cast_354_wire_constant when (BITSEL_u8_u1_352_wire(0) /=  '0') else type_cast_356_wire_constant;
    -- flow-through select operator MUX_367_inst
    IMA19_368 <= type_cast_364_wire_constant when (BITSEL_u8_u1_362_wire(0) /=  '0') else type_cast_366_wire_constant;
    -- flow-through select operator MUX_377_inst
    IMA20_378 <= type_cast_374_wire_constant when (BITSEL_u8_u1_372_wire(0) /=  '0') else type_cast_376_wire_constant;
    -- flow-through select operator MUX_387_inst
    IMA21_388 <= type_cast_384_wire_constant when (BITSEL_u8_u1_382_wire(0) /=  '0') else type_cast_386_wire_constant;
    -- flow-through select operator MUX_397_inst
    IMA22_398 <= type_cast_394_wire_constant when (BITSEL_u8_u1_392_wire(0) /=  '0') else type_cast_396_wire_constant;
    -- flow-through select operator MUX_407_inst
    IMA23_408 <= type_cast_404_wire_constant when (BITSEL_u8_u1_402_wire(0) /=  '0') else type_cast_406_wire_constant;
    -- flow-through select operator MUX_417_inst
    IMA24_418 <= type_cast_414_wire_constant when (BITSEL_u8_u1_412_wire(0) /=  '0') else type_cast_416_wire_constant;
    -- flow-through select operator MUX_427_inst
    IMA25_428 <= type_cast_424_wire_constant when (BITSEL_u8_u1_422_wire(0) /=  '0') else type_cast_426_wire_constant;
    -- flow-through select operator MUX_437_inst
    IMA26_438 <= type_cast_434_wire_constant when (BITSEL_u8_u1_432_wire(0) /=  '0') else type_cast_436_wire_constant;
    -- flow-through select operator MUX_447_inst
    IMA27_448 <= type_cast_444_wire_constant when (BITSEL_u8_u1_442_wire(0) /=  '0') else type_cast_446_wire_constant;
    -- flow-through select operator MUX_457_inst
    IMA28_458 <= type_cast_454_wire_constant when (BITSEL_u8_u1_452_wire(0) /=  '0') else type_cast_456_wire_constant;
    -- flow-through select operator MUX_467_inst
    IMA29_468 <= type_cast_464_wire_constant when (BITSEL_u8_u1_462_wire(0) /=  '0') else type_cast_466_wire_constant;
    -- flow-through select operator MUX_477_inst
    IMA30_478 <= type_cast_474_wire_constant when (BITSEL_u8_u1_472_wire(0) /=  '0') else type_cast_476_wire_constant;
    -- flow-through select operator MUX_487_inst
    IMA31_488 <= type_cast_484_wire_constant when (BITSEL_u8_u1_482_wire(0) /=  '0') else type_cast_486_wire_constant;
    -- flow-through select operator MUX_497_inst
    IMA32_498 <= type_cast_494_wire_constant when (BITSEL_u8_u1_492_wire(0) /=  '0') else type_cast_496_wire_constant;
    -- flow-through select operator MUX_507_inst
    IMA33_508 <= type_cast_504_wire_constant when (BITSEL_u8_u1_502_wire(0) /=  '0') else type_cast_506_wire_constant;
    -- flow-through select operator MUX_517_inst
    IMA34_518 <= type_cast_514_wire_constant when (BITSEL_u8_u1_512_wire(0) /=  '0') else type_cast_516_wire_constant;
    -- flow-through select operator MUX_527_inst
    IMA35_528 <= type_cast_524_wire_constant when (BITSEL_u8_u1_522_wire(0) /=  '0') else type_cast_526_wire_constant;
    -- flow-through select operator MUX_537_inst
    IMA36_538 <= type_cast_534_wire_constant when (BITSEL_u8_u1_532_wire(0) /=  '0') else type_cast_536_wire_constant;
    -- flow-through select operator MUX_547_inst
    IMA37_548 <= type_cast_544_wire_constant when (BITSEL_u8_u1_542_wire(0) /=  '0') else type_cast_546_wire_constant;
    -- flow-through select operator MUX_557_inst
    IMA38_558 <= type_cast_554_wire_constant when (BITSEL_u8_u1_552_wire(0) /=  '0') else type_cast_556_wire_constant;
    -- flow-through select operator MUX_567_inst
    IMA39_568 <= type_cast_564_wire_constant when (BITSEL_u8_u1_562_wire(0) /=  '0') else type_cast_566_wire_constant;
    -- flow-through select operator MUX_577_inst
    IMA40_578 <= type_cast_574_wire_constant when (BITSEL_u8_u1_572_wire(0) /=  '0') else type_cast_576_wire_constant;
    -- flow-through select operator MUX_587_inst
    IMA41_588 <= type_cast_584_wire_constant when (BITSEL_u8_u1_582_wire(0) /=  '0') else type_cast_586_wire_constant;
    -- flow-through select operator MUX_597_inst
    IMA42_598 <= type_cast_594_wire_constant when (BITSEL_u8_u1_592_wire(0) /=  '0') else type_cast_596_wire_constant;
    -- flow-through select operator MUX_607_inst
    IMA43_608 <= type_cast_604_wire_constant when (BITSEL_u8_u1_602_wire(0) /=  '0') else type_cast_606_wire_constant;
    -- flow-through select operator MUX_617_inst
    IMA44_618 <= type_cast_614_wire_constant when (BITSEL_u8_u1_612_wire(0) /=  '0') else type_cast_616_wire_constant;
    -- flow-through select operator MUX_627_inst
    IMA45_628 <= type_cast_624_wire_constant when (BITSEL_u8_u1_622_wire(0) /=  '0') else type_cast_626_wire_constant;
    -- flow-through select operator MUX_637_inst
    IMA46_638 <= type_cast_634_wire_constant when (BITSEL_u8_u1_632_wire(0) /=  '0') else type_cast_636_wire_constant;
    -- flow-through select operator MUX_647_inst
    IMA47_648 <= type_cast_644_wire_constant when (BITSEL_u8_u1_642_wire(0) /=  '0') else type_cast_646_wire_constant;
    -- flow-through select operator MUX_657_inst
    IMA48_658 <= type_cast_654_wire_constant when (BITSEL_u8_u1_652_wire(0) /=  '0') else type_cast_656_wire_constant;
    -- flow-through select operator MUX_667_inst
    IMA49_668 <= type_cast_664_wire_constant when (BITSEL_u8_u1_662_wire(0) /=  '0') else type_cast_666_wire_constant;
    -- flow-through select operator MUX_677_inst
    IMA50_678 <= type_cast_674_wire_constant when (BITSEL_u8_u1_672_wire(0) /=  '0') else type_cast_676_wire_constant;
    -- flow-through select operator MUX_687_inst
    IMA51_688 <= type_cast_684_wire_constant when (BITSEL_u8_u1_682_wire(0) /=  '0') else type_cast_686_wire_constant;
    -- flow-through select operator MUX_697_inst
    IMA52_698 <= type_cast_694_wire_constant when (BITSEL_u8_u1_692_wire(0) /=  '0') else type_cast_696_wire_constant;
    -- flow-through select operator MUX_707_inst
    IMA53_708 <= type_cast_704_wire_constant when (BITSEL_u8_u1_702_wire(0) /=  '0') else type_cast_706_wire_constant;
    -- flow-through select operator MUX_717_inst
    IMA54_718 <= type_cast_714_wire_constant when (BITSEL_u8_u1_712_wire(0) /=  '0') else type_cast_716_wire_constant;
    -- flow-through select operator MUX_727_inst
    IMA55_728 <= type_cast_724_wire_constant when (BITSEL_u8_u1_722_wire(0) /=  '0') else type_cast_726_wire_constant;
    -- flow-through select operator MUX_737_inst
    IMA56_738 <= type_cast_734_wire_constant when (BITSEL_u8_u1_732_wire(0) /=  '0') else type_cast_736_wire_constant;
    -- flow-through select operator MUX_747_inst
    IMA57_748 <= type_cast_744_wire_constant when (BITSEL_u8_u1_742_wire(0) /=  '0') else type_cast_746_wire_constant;
    -- flow-through select operator MUX_757_inst
    IMA58_758 <= type_cast_754_wire_constant when (BITSEL_u8_u1_752_wire(0) /=  '0') else type_cast_756_wire_constant;
    -- flow-through select operator MUX_767_inst
    IMA59_768 <= type_cast_764_wire_constant when (BITSEL_u8_u1_762_wire(0) /=  '0') else type_cast_766_wire_constant;
    -- flow-through select operator MUX_777_inst
    IMA60_778 <= type_cast_774_wire_constant when (BITSEL_u8_u1_772_wire(0) /=  '0') else type_cast_776_wire_constant;
    -- flow-through select operator MUX_787_inst
    IMA61_788 <= type_cast_784_wire_constant when (BITSEL_u8_u1_782_wire(0) /=  '0') else type_cast_786_wire_constant;
    -- flow-through select operator MUX_797_inst
    IMA62_798 <= type_cast_794_wire_constant when (BITSEL_u8_u1_792_wire(0) /=  '0') else type_cast_796_wire_constant;
    -- flow-through select operator MUX_807_inst
    IMA63_808 <= type_cast_804_wire_constant when (BITSEL_u8_u1_802_wire(0) /=  '0') else type_cast_806_wire_constant;
    -- flow-through select operator MUX_817_inst
    IMA64_818 <= type_cast_814_wire_constant when (BITSEL_u8_u1_812_wire(0) /=  '0') else type_cast_816_wire_constant;
    -- flow-through select operator MUX_827_inst
    IMA65_828 <= type_cast_824_wire_constant when (BITSEL_u8_u1_822_wire(0) /=  '0') else type_cast_826_wire_constant;
    -- flow-through select operator MUX_837_inst
    IMA66_838 <= type_cast_834_wire_constant when (BITSEL_u8_u1_832_wire(0) /=  '0') else type_cast_836_wire_constant;
    -- flow-through select operator MUX_847_inst
    IMA67_848 <= type_cast_844_wire_constant when (BITSEL_u8_u1_842_wire(0) /=  '0') else type_cast_846_wire_constant;
    -- flow-through select operator MUX_857_inst
    IMA68_858 <= type_cast_854_wire_constant when (BITSEL_u8_u1_852_wire(0) /=  '0') else type_cast_856_wire_constant;
    -- flow-through select operator MUX_867_inst
    IMA69_868 <= type_cast_864_wire_constant when (BITSEL_u8_u1_862_wire(0) /=  '0') else type_cast_866_wire_constant;
    -- flow-through select operator MUX_877_inst
    IMA70_878 <= type_cast_874_wire_constant when (BITSEL_u8_u1_872_wire(0) /=  '0') else type_cast_876_wire_constant;
    -- flow-through select operator MUX_887_inst
    IMA71_888 <= type_cast_884_wire_constant when (BITSEL_u8_u1_882_wire(0) /=  '0') else type_cast_886_wire_constant;
    -- flow-through select operator MUX_897_inst
    IMA72_898 <= type_cast_894_wire_constant when (BITSEL_u8_u1_892_wire(0) /=  '0') else type_cast_896_wire_constant;
    -- flow-through select operator MUX_907_inst
    IMA73_908 <= type_cast_904_wire_constant when (BITSEL_u8_u1_902_wire(0) /=  '0') else type_cast_906_wire_constant;
    -- flow-through select operator MUX_917_inst
    IMA74_918 <= type_cast_914_wire_constant when (BITSEL_u8_u1_912_wire(0) /=  '0') else type_cast_916_wire_constant;
    -- flow-through select operator MUX_927_inst
    IMA75_928 <= type_cast_924_wire_constant when (BITSEL_u8_u1_922_wire(0) /=  '0') else type_cast_926_wire_constant;
    -- flow-through select operator MUX_937_inst
    IMA76_938 <= type_cast_934_wire_constant when (BITSEL_u8_u1_932_wire(0) /=  '0') else type_cast_936_wire_constant;
    -- flow-through select operator MUX_947_inst
    IMA77_948 <= type_cast_944_wire_constant when (BITSEL_u8_u1_942_wire(0) /=  '0') else type_cast_946_wire_constant;
    -- flow-through select operator MUX_957_inst
    IMA78_958 <= type_cast_954_wire_constant when (BITSEL_u8_u1_952_wire(0) /=  '0') else type_cast_956_wire_constant;
    -- flow-through select operator MUX_967_inst
    IMA79_968 <= type_cast_964_wire_constant when (BITSEL_u8_u1_962_wire(0) /=  '0') else type_cast_966_wire_constant;
    -- flow-through select operator MUX_977_inst
    IMA80_978 <= type_cast_974_wire_constant when (BITSEL_u8_u1_972_wire(0) /=  '0') else type_cast_976_wire_constant;
    -- flow-through select operator MUX_987_inst
    IMA81_988 <= type_cast_984_wire_constant when (BITSEL_u8_u1_982_wire(0) /=  '0') else type_cast_986_wire_constant;
    -- flow-through select operator MUX_997_inst
    IMA82_998 <= type_cast_994_wire_constant when (BITSEL_u8_u1_992_wire(0) /=  '0') else type_cast_996_wire_constant;
    -- binary operator BITSEL_u8_u1_1002_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1001_wire_constant, tmp_var);
      BITSEL_u8_u1_1002_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1012_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1011_wire_constant, tmp_var);
      BITSEL_u8_u1_1012_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1022_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1021_wire_constant, tmp_var);
      BITSEL_u8_u1_1022_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1032_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1031_wire_constant, tmp_var);
      BITSEL_u8_u1_1032_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1042_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1041_wire_constant, tmp_var);
      BITSEL_u8_u1_1042_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1052_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1051_wire_constant, tmp_var);
      BITSEL_u8_u1_1052_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1062_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1061_wire_constant, tmp_var);
      BITSEL_u8_u1_1062_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1072_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1071_wire_constant, tmp_var);
      BITSEL_u8_u1_1072_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1082_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1081_wire_constant, tmp_var);
      BITSEL_u8_u1_1082_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1092_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1091_wire_constant, tmp_var);
      BITSEL_u8_u1_1092_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1102_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1101_wire_constant, tmp_var);
      BITSEL_u8_u1_1102_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1112_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1111_wire_constant, tmp_var);
      BITSEL_u8_u1_1112_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1122_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1121_wire_constant, tmp_var);
      BITSEL_u8_u1_1122_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1132_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1131_wire_constant, tmp_var);
      BITSEL_u8_u1_1132_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1142_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1141_wire_constant, tmp_var);
      BITSEL_u8_u1_1142_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1152_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1151_wire_constant, tmp_var);
      BITSEL_u8_u1_1152_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1162_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1161_wire_constant, tmp_var);
      BITSEL_u8_u1_1162_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1172_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1171_wire_constant, tmp_var);
      BITSEL_u8_u1_1172_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1182_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1181_wire_constant, tmp_var);
      BITSEL_u8_u1_1182_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1192_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1191_wire_constant, tmp_var);
      BITSEL_u8_u1_1192_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1202_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1201_wire_constant, tmp_var);
      BITSEL_u8_u1_1202_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1212_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1211_wire_constant, tmp_var);
      BITSEL_u8_u1_1212_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1222_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1221_wire_constant, tmp_var);
      BITSEL_u8_u1_1222_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1232_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1231_wire_constant, tmp_var);
      BITSEL_u8_u1_1232_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1242_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1241_wire_constant, tmp_var);
      BITSEL_u8_u1_1242_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1252_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1251_wire_constant, tmp_var);
      BITSEL_u8_u1_1252_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1262_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1261_wire_constant, tmp_var);
      BITSEL_u8_u1_1262_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1272_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1271_wire_constant, tmp_var);
      BITSEL_u8_u1_1272_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1282_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1281_wire_constant, tmp_var);
      BITSEL_u8_u1_1282_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1292_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1291_wire_constant, tmp_var);
      BITSEL_u8_u1_1292_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1302_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1301_wire_constant, tmp_var);
      BITSEL_u8_u1_1302_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1312_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1311_wire_constant, tmp_var);
      BITSEL_u8_u1_1312_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1322_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1321_wire_constant, tmp_var);
      BITSEL_u8_u1_1322_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1332_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1331_wire_constant, tmp_var);
      BITSEL_u8_u1_1332_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1342_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1341_wire_constant, tmp_var);
      BITSEL_u8_u1_1342_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1352_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1351_wire_constant, tmp_var);
      BITSEL_u8_u1_1352_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1362_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1361_wire_constant, tmp_var);
      BITSEL_u8_u1_1362_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1372_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1371_wire_constant, tmp_var);
      BITSEL_u8_u1_1372_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1382_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1381_wire_constant, tmp_var);
      BITSEL_u8_u1_1382_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1392_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1391_wire_constant, tmp_var);
      BITSEL_u8_u1_1392_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1402_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1401_wire_constant, tmp_var);
      BITSEL_u8_u1_1402_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1412_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1411_wire_constant, tmp_var);
      BITSEL_u8_u1_1412_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1422_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1421_wire_constant, tmp_var);
      BITSEL_u8_u1_1422_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1432_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1431_wire_constant, tmp_var);
      BITSEL_u8_u1_1432_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1442_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1441_wire_constant, tmp_var);
      BITSEL_u8_u1_1442_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1452_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1451_wire_constant, tmp_var);
      BITSEL_u8_u1_1452_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1460_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1459_wire_constant, tmp_var);
      BITSEL_u8_u1_1460_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1468_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1467_wire_constant, tmp_var);
      BITSEL_u8_u1_1468_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1476_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1475_wire_constant, tmp_var);
      BITSEL_u8_u1_1476_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1484_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1483_wire_constant, tmp_var);
      BITSEL_u8_u1_1484_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1492_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1491_wire_constant, tmp_var);
      BITSEL_u8_u1_1492_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1500_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1499_wire_constant, tmp_var);
      BITSEL_u8_u1_1500_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1508_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1507_wire_constant, tmp_var);
      BITSEL_u8_u1_1508_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1516_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1515_wire_constant, tmp_var);
      BITSEL_u8_u1_1516_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1524_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1523_wire_constant, tmp_var);
      BITSEL_u8_u1_1524_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1532_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1531_wire_constant, tmp_var);
      BITSEL_u8_u1_1532_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1540_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1539_wire_constant, tmp_var);
      BITSEL_u8_u1_1540_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1548_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1547_wire_constant, tmp_var);
      BITSEL_u8_u1_1548_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1556_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1555_wire_constant, tmp_var);
      BITSEL_u8_u1_1556_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1564_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1563_wire_constant, tmp_var);
      BITSEL_u8_u1_1564_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1572_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1571_wire_constant, tmp_var);
      BITSEL_u8_u1_1572_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1580_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1579_wire_constant, tmp_var);
      BITSEL_u8_u1_1580_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1588_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1587_wire_constant, tmp_var);
      BITSEL_u8_u1_1588_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1596_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1595_wire_constant, tmp_var);
      BITSEL_u8_u1_1596_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1604_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1603_wire_constant, tmp_var);
      BITSEL_u8_u1_1604_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1612_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1611_wire_constant, tmp_var);
      BITSEL_u8_u1_1612_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1620_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1619_wire_constant, tmp_var);
      BITSEL_u8_u1_1620_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1628_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1627_wire_constant, tmp_var);
      BITSEL_u8_u1_1628_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1636_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1635_wire_constant, tmp_var);
      BITSEL_u8_u1_1636_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1644_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1643_wire_constant, tmp_var);
      BITSEL_u8_u1_1644_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1652_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1651_wire_constant, tmp_var);
      BITSEL_u8_u1_1652_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1660_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1659_wire_constant, tmp_var);
      BITSEL_u8_u1_1660_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1668_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1667_wire_constant, tmp_var);
      BITSEL_u8_u1_1668_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1676_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1675_wire_constant, tmp_var);
      BITSEL_u8_u1_1676_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1684_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1683_wire_constant, tmp_var);
      BITSEL_u8_u1_1684_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1692_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1691_wire_constant, tmp_var);
      BITSEL_u8_u1_1692_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1700_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1699_wire_constant, tmp_var);
      BITSEL_u8_u1_1700_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1708_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1707_wire_constant, tmp_var);
      BITSEL_u8_u1_1708_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1716_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1715_wire_constant, tmp_var);
      BITSEL_u8_u1_1716_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1724_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1723_wire_constant, tmp_var);
      BITSEL_u8_u1_1724_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_172_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_171_wire_constant, tmp_var);
      BITSEL_u8_u1_172_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1732_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1731_wire_constant, tmp_var);
      BITSEL_u8_u1_1732_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1740_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1739_wire_constant, tmp_var);
      BITSEL_u8_u1_1740_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1748_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1747_wire_constant, tmp_var);
      BITSEL_u8_u1_1748_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1756_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1755_wire_constant, tmp_var);
      BITSEL_u8_u1_1756_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1764_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1763_wire_constant, tmp_var);
      BITSEL_u8_u1_1764_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1772_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1771_wire_constant, tmp_var);
      BITSEL_u8_u1_1772_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1780_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1779_wire_constant, tmp_var);
      BITSEL_u8_u1_1780_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1788_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1787_wire_constant, tmp_var);
      BITSEL_u8_u1_1788_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1796_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1795_wire_constant, tmp_var);
      BITSEL_u8_u1_1796_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1804_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1803_wire_constant, tmp_var);
      BITSEL_u8_u1_1804_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1812_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1811_wire_constant, tmp_var);
      BITSEL_u8_u1_1812_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1820_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1819_wire_constant, tmp_var);
      BITSEL_u8_u1_1820_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1828_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1827_wire_constant, tmp_var);
      BITSEL_u8_u1_1828_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_182_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_181_wire_constant, tmp_var);
      BITSEL_u8_u1_182_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1836_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1835_wire_constant, tmp_var);
      BITSEL_u8_u1_1836_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1844_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1843_wire_constant, tmp_var);
      BITSEL_u8_u1_1844_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1852_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1851_wire_constant, tmp_var);
      BITSEL_u8_u1_1852_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1860_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1859_wire_constant, tmp_var);
      BITSEL_u8_u1_1860_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1868_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1867_wire_constant, tmp_var);
      BITSEL_u8_u1_1868_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1876_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1875_wire_constant, tmp_var);
      BITSEL_u8_u1_1876_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1884_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1883_wire_constant, tmp_var);
      BITSEL_u8_u1_1884_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1892_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1891_wire_constant, tmp_var);
      BITSEL_u8_u1_1892_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1900_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1899_wire_constant, tmp_var);
      BITSEL_u8_u1_1900_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1908_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1907_wire_constant, tmp_var);
      BITSEL_u8_u1_1908_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1916_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1915_wire_constant, tmp_var);
      BITSEL_u8_u1_1916_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1924_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1923_wire_constant, tmp_var);
      BITSEL_u8_u1_1924_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_192_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_191_wire_constant, tmp_var);
      BITSEL_u8_u1_192_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1932_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1931_wire_constant, tmp_var);
      BITSEL_u8_u1_1932_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1940_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1939_wire_constant, tmp_var);
      BITSEL_u8_u1_1940_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1948_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1947_wire_constant, tmp_var);
      BITSEL_u8_u1_1948_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1956_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1955_wire_constant, tmp_var);
      BITSEL_u8_u1_1956_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1964_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1963_wire_constant, tmp_var);
      BITSEL_u8_u1_1964_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1972_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1971_wire_constant, tmp_var);
      BITSEL_u8_u1_1972_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1980_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1979_wire_constant, tmp_var);
      BITSEL_u8_u1_1980_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1988_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1987_wire_constant, tmp_var);
      BITSEL_u8_u1_1988_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1996_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_1995_wire_constant, tmp_var);
      BITSEL_u8_u1_1996_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2004_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2003_wire_constant, tmp_var);
      BITSEL_u8_u1_2004_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2012_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2011_wire_constant, tmp_var);
      BITSEL_u8_u1_2012_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2020_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2019_wire_constant, tmp_var);
      BITSEL_u8_u1_2020_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2028_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2027_wire_constant, tmp_var);
      BITSEL_u8_u1_2028_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_202_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_201_wire_constant, tmp_var);
      BITSEL_u8_u1_202_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2036_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2035_wire_constant, tmp_var);
      BITSEL_u8_u1_2036_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2044_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2043_wire_constant, tmp_var);
      BITSEL_u8_u1_2044_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2052_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2051_wire_constant, tmp_var);
      BITSEL_u8_u1_2052_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2060_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2059_wire_constant, tmp_var);
      BITSEL_u8_u1_2060_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2068_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2067_wire_constant, tmp_var);
      BITSEL_u8_u1_2068_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2076_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2075_wire_constant, tmp_var);
      BITSEL_u8_u1_2076_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2084_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2083_wire_constant, tmp_var);
      BITSEL_u8_u1_2084_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2092_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2091_wire_constant, tmp_var);
      BITSEL_u8_u1_2092_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2100_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2099_wire_constant, tmp_var);
      BITSEL_u8_u1_2100_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2108_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2107_wire_constant, tmp_var);
      BITSEL_u8_u1_2108_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2116_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2115_wire_constant, tmp_var);
      BITSEL_u8_u1_2116_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2124_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2123_wire_constant, tmp_var);
      BITSEL_u8_u1_2124_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_212_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_211_wire_constant, tmp_var);
      BITSEL_u8_u1_212_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2132_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2131_wire_constant, tmp_var);
      BITSEL_u8_u1_2132_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2140_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2139_wire_constant, tmp_var);
      BITSEL_u8_u1_2140_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2148_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2147_wire_constant, tmp_var);
      BITSEL_u8_u1_2148_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2156_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2155_wire_constant, tmp_var);
      BITSEL_u8_u1_2156_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2164_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2163_wire_constant, tmp_var);
      BITSEL_u8_u1_2164_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2172_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2171_wire_constant, tmp_var);
      BITSEL_u8_u1_2172_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2180_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2179_wire_constant, tmp_var);
      BITSEL_u8_u1_2180_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2188_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2187_wire_constant, tmp_var);
      BITSEL_u8_u1_2188_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2196_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2195_wire_constant, tmp_var);
      BITSEL_u8_u1_2196_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2204_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2203_wire_constant, tmp_var);
      BITSEL_u8_u1_2204_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2212_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2211_wire_constant, tmp_var);
      BITSEL_u8_u1_2212_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2220_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2219_wire_constant, tmp_var);
      BITSEL_u8_u1_2220_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2228_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2227_wire_constant, tmp_var);
      BITSEL_u8_u1_2228_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_222_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_221_wire_constant, tmp_var);
      BITSEL_u8_u1_222_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2236_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2235_wire_constant, tmp_var);
      BITSEL_u8_u1_2236_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2244_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2243_wire_constant, tmp_var);
      BITSEL_u8_u1_2244_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2252_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2251_wire_constant, tmp_var);
      BITSEL_u8_u1_2252_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2260_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2259_wire_constant, tmp_var);
      BITSEL_u8_u1_2260_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2268_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2267_wire_constant, tmp_var);
      BITSEL_u8_u1_2268_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2276_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2275_wire_constant, tmp_var);
      BITSEL_u8_u1_2276_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2284_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2283_wire_constant, tmp_var);
      BITSEL_u8_u1_2284_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2292_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2291_wire_constant, tmp_var);
      BITSEL_u8_u1_2292_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2300_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2299_wire_constant, tmp_var);
      BITSEL_u8_u1_2300_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2308_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2307_wire_constant, tmp_var);
      BITSEL_u8_u1_2308_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2316_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2315_wire_constant, tmp_var);
      BITSEL_u8_u1_2316_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2324_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2323_wire_constant, tmp_var);
      BITSEL_u8_u1_2324_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_232_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_231_wire_constant, tmp_var);
      BITSEL_u8_u1_232_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2332_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2331_wire_constant, tmp_var);
      BITSEL_u8_u1_2332_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2340_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2339_wire_constant, tmp_var);
      BITSEL_u8_u1_2340_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2348_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2347_wire_constant, tmp_var);
      BITSEL_u8_u1_2348_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2356_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2355_wire_constant, tmp_var);
      BITSEL_u8_u1_2356_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2364_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2363_wire_constant, tmp_var);
      BITSEL_u8_u1_2364_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2372_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2371_wire_constant, tmp_var);
      BITSEL_u8_u1_2372_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2380_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2379_wire_constant, tmp_var);
      BITSEL_u8_u1_2380_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2388_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2387_wire_constant, tmp_var);
      BITSEL_u8_u1_2388_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2396_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2395_wire_constant, tmp_var);
      BITSEL_u8_u1_2396_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2404_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2403_wire_constant, tmp_var);
      BITSEL_u8_u1_2404_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2412_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2411_wire_constant, tmp_var);
      BITSEL_u8_u1_2412_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2420_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2419_wire_constant, tmp_var);
      BITSEL_u8_u1_2420_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2428_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2427_wire_constant, tmp_var);
      BITSEL_u8_u1_2428_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_242_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_241_wire_constant, tmp_var);
      BITSEL_u8_u1_242_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2436_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2435_wire_constant, tmp_var);
      BITSEL_u8_u1_2436_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2444_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2443_wire_constant, tmp_var);
      BITSEL_u8_u1_2444_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2452_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2451_wire_constant, tmp_var);
      BITSEL_u8_u1_2452_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2460_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2459_wire_constant, tmp_var);
      BITSEL_u8_u1_2460_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_252_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_251_wire_constant, tmp_var);
      BITSEL_u8_u1_252_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_262_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_261_wire_constant, tmp_var);
      BITSEL_u8_u1_262_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_272_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_271_wire_constant, tmp_var);
      BITSEL_u8_u1_272_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_282_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_281_wire_constant, tmp_var);
      BITSEL_u8_u1_282_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_292_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_291_wire_constant, tmp_var);
      BITSEL_u8_u1_292_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_302_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_301_wire_constant, tmp_var);
      BITSEL_u8_u1_302_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_312_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_311_wire_constant, tmp_var);
      BITSEL_u8_u1_312_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_322_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_321_wire_constant, tmp_var);
      BITSEL_u8_u1_322_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_332_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_331_wire_constant, tmp_var);
      BITSEL_u8_u1_332_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_342_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_341_wire_constant, tmp_var);
      BITSEL_u8_u1_342_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_352_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_351_wire_constant, tmp_var);
      BITSEL_u8_u1_352_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_362_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_361_wire_constant, tmp_var);
      BITSEL_u8_u1_362_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_372_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_371_wire_constant, tmp_var);
      BITSEL_u8_u1_372_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_382_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_381_wire_constant, tmp_var);
      BITSEL_u8_u1_382_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_392_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_391_wire_constant, tmp_var);
      BITSEL_u8_u1_392_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_402_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_401_wire_constant, tmp_var);
      BITSEL_u8_u1_402_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_412_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_411_wire_constant, tmp_var);
      BITSEL_u8_u1_412_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_422_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_421_wire_constant, tmp_var);
      BITSEL_u8_u1_422_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_432_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_431_wire_constant, tmp_var);
      BITSEL_u8_u1_432_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_442_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_441_wire_constant, tmp_var);
      BITSEL_u8_u1_442_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_452_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_451_wire_constant, tmp_var);
      BITSEL_u8_u1_452_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_462_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_461_wire_constant, tmp_var);
      BITSEL_u8_u1_462_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_472_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_471_wire_constant, tmp_var);
      BITSEL_u8_u1_472_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_482_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_481_wire_constant, tmp_var);
      BITSEL_u8_u1_482_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_492_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_491_wire_constant, tmp_var);
      BITSEL_u8_u1_492_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_502_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_501_wire_constant, tmp_var);
      BITSEL_u8_u1_502_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_512_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_511_wire_constant, tmp_var);
      BITSEL_u8_u1_512_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_522_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_521_wire_constant, tmp_var);
      BITSEL_u8_u1_522_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_532_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_531_wire_constant, tmp_var);
      BITSEL_u8_u1_532_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_542_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_541_wire_constant, tmp_var);
      BITSEL_u8_u1_542_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_552_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_551_wire_constant, tmp_var);
      BITSEL_u8_u1_552_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_562_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_561_wire_constant, tmp_var);
      BITSEL_u8_u1_562_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_572_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_571_wire_constant, tmp_var);
      BITSEL_u8_u1_572_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_582_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_581_wire_constant, tmp_var);
      BITSEL_u8_u1_582_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_592_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_591_wire_constant, tmp_var);
      BITSEL_u8_u1_592_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_602_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_601_wire_constant, tmp_var);
      BITSEL_u8_u1_602_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_612_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_611_wire_constant, tmp_var);
      BITSEL_u8_u1_612_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_622_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_621_wire_constant, tmp_var);
      BITSEL_u8_u1_622_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_632_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_631_wire_constant, tmp_var);
      BITSEL_u8_u1_632_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_642_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_641_wire_constant, tmp_var);
      BITSEL_u8_u1_642_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_652_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_651_wire_constant, tmp_var);
      BITSEL_u8_u1_652_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_662_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_661_wire_constant, tmp_var);
      BITSEL_u8_u1_662_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_672_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_671_wire_constant, tmp_var);
      BITSEL_u8_u1_672_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_682_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_681_wire_constant, tmp_var);
      BITSEL_u8_u1_682_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_692_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_691_wire_constant, tmp_var);
      BITSEL_u8_u1_692_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_702_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_701_wire_constant, tmp_var);
      BITSEL_u8_u1_702_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_712_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_711_wire_constant, tmp_var);
      BITSEL_u8_u1_712_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_722_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_721_wire_constant, tmp_var);
      BITSEL_u8_u1_722_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_732_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_731_wire_constant, tmp_var);
      BITSEL_u8_u1_732_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_742_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_741_wire_constant, tmp_var);
      BITSEL_u8_u1_742_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_752_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_751_wire_constant, tmp_var);
      BITSEL_u8_u1_752_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_762_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_761_wire_constant, tmp_var);
      BITSEL_u8_u1_762_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_772_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_771_wire_constant, tmp_var);
      BITSEL_u8_u1_772_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_782_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_781_wire_constant, tmp_var);
      BITSEL_u8_u1_782_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_792_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_791_wire_constant, tmp_var);
      BITSEL_u8_u1_792_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_802_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_801_wire_constant, tmp_var);
      BITSEL_u8_u1_802_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_812_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_811_wire_constant, tmp_var);
      BITSEL_u8_u1_812_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_822_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_821_wire_constant, tmp_var);
      BITSEL_u8_u1_822_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_832_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_831_wire_constant, tmp_var);
      BITSEL_u8_u1_832_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_842_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_841_wire_constant, tmp_var);
      BITSEL_u8_u1_842_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_852_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_851_wire_constant, tmp_var);
      BITSEL_u8_u1_852_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_862_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_861_wire_constant, tmp_var);
      BITSEL_u8_u1_862_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_872_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_871_wire_constant, tmp_var);
      BITSEL_u8_u1_872_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_882_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_881_wire_constant, tmp_var);
      BITSEL_u8_u1_882_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_892_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_891_wire_constant, tmp_var);
      BITSEL_u8_u1_892_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_902_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_901_wire_constant, tmp_var);
      BITSEL_u8_u1_902_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_912_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_911_wire_constant, tmp_var);
      BITSEL_u8_u1_912_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_922_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_921_wire_constant, tmp_var);
      BITSEL_u8_u1_922_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_932_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_931_wire_constant, tmp_var);
      BITSEL_u8_u1_932_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_942_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_941_wire_constant, tmp_var);
      BITSEL_u8_u1_942_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_952_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_951_wire_constant, tmp_var);
      BITSEL_u8_u1_952_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_962_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_961_wire_constant, tmp_var);
      BITSEL_u8_u1_962_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_972_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_971_wire_constant, tmp_var);
      BITSEL_u8_u1_972_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_982_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_981_wire_constant, tmp_var);
      BITSEL_u8_u1_982_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_992_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_991_wire_constant, tmp_var);
      BITSEL_u8_u1_992_wire <= tmp_var; -- 
    end process;
    -- 
  end Block; -- data_path
  -- 
end Inv_Sbox_1_Volatile_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library work;
use work.ahir_system_global_package.all;
entity Inv_Sbox_2_Volatile is -- 
  port ( -- 
    s_in : in  std_logic_vector(7 downto 0);
    s_out : out  std_logic_vector(7 downto 0)-- 
  );
  -- 
end entity Inv_Sbox_2_Volatile;
architecture Inv_Sbox_2_Volatile_arch of Inv_Sbox_2_Volatile is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector(8-1 downto 0);
  signal default_zero_sig: std_logic;
  -- input port buffer signals
  signal s_in_buffer :  std_logic_vector(7 downto 0);
  -- output port buffer signals
  signal s_out_buffer :  std_logic_vector(7 downto 0);
  -- volatile/operator module components. 
  -- 
begin --  
  -- input handling ------------------------------------------------
  s_in_buffer <= s_in;
  -- output handling  -------------------------------------------------------
  s_out <= s_out_buffer;
  -- the control path --------------------------------------------------
  default_zero_sig <= '0';
  -- volatile module, no control path
  -- the data path
  data_path: Block -- 
    signal BITSEL_u8_u1_2472_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2482_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2492_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2502_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2512_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2522_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2532_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2542_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2552_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2562_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2572_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2582_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2592_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2602_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2612_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2622_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2632_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2642_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2652_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2662_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2672_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2682_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2692_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2702_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2712_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2722_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2732_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2742_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2752_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2762_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2772_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2782_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2792_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2802_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2812_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2822_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2832_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2842_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2852_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2862_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2872_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2882_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2892_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2902_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2912_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2922_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2932_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2942_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2952_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2962_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2972_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2982_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_2992_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3002_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3012_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3022_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3032_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3042_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3052_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3062_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3072_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3082_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3092_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3102_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3112_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3122_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3132_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3142_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3152_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3162_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3172_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3182_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3192_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3202_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3212_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3222_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3232_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3242_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3252_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3262_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3272_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3282_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3292_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3302_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3312_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3322_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3332_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3342_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3352_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3362_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3372_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3382_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3392_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3402_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3412_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3422_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3432_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3442_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3452_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3462_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3472_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3482_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3492_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3502_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3512_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3522_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3532_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3542_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3552_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3562_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3572_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3582_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3592_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3602_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3612_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3622_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3632_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3642_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3652_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3662_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3672_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3682_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3692_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3702_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3712_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3722_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3732_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3742_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3752_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3760_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3768_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3776_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3784_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3792_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3800_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3808_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3816_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3824_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3832_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3840_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3848_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3856_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3864_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3872_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3880_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3888_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3896_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3904_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3912_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3920_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3928_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3936_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3944_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3952_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3960_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3968_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3976_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3984_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_3992_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4000_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4008_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4016_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4024_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4032_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4040_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4048_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4056_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4064_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4072_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4080_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4088_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4096_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4104_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4112_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4120_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4128_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4136_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4144_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4152_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4160_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4168_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4176_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4184_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4192_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4200_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4208_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4216_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4224_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4232_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4240_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4248_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4256_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4264_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4272_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4280_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4288_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4296_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4304_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4312_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4320_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4328_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4336_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4344_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4352_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4360_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4368_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4376_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4384_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4392_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4400_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4408_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4416_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4424_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4432_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4440_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4448_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4456_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4464_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4472_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4480_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4488_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4496_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4504_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4512_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4520_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4528_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4536_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4544_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4552_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4560_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4568_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4576_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4584_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4592_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4600_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4608_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4616_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4624_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4632_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4640_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4648_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4656_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4664_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4672_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4680_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4688_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4696_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4704_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4712_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4720_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4728_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4736_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4744_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4752_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4760_wire : std_logic_vector(0 downto 0);
    signal IMA0_2478 : std_logic_vector(7 downto 0);
    signal IMA100_3478 : std_logic_vector(7 downto 0);
    signal IMA101_3488 : std_logic_vector(7 downto 0);
    signal IMA102_3498 : std_logic_vector(7 downto 0);
    signal IMA103_3508 : std_logic_vector(7 downto 0);
    signal IMA104_3518 : std_logic_vector(7 downto 0);
    signal IMA105_3528 : std_logic_vector(7 downto 0);
    signal IMA106_3538 : std_logic_vector(7 downto 0);
    signal IMA107_3548 : std_logic_vector(7 downto 0);
    signal IMA108_3558 : std_logic_vector(7 downto 0);
    signal IMA109_3568 : std_logic_vector(7 downto 0);
    signal IMA10_2578 : std_logic_vector(7 downto 0);
    signal IMA110_3578 : std_logic_vector(7 downto 0);
    signal IMA111_3588 : std_logic_vector(7 downto 0);
    signal IMA112_3598 : std_logic_vector(7 downto 0);
    signal IMA113_3608 : std_logic_vector(7 downto 0);
    signal IMA114_3618 : std_logic_vector(7 downto 0);
    signal IMA115_3628 : std_logic_vector(7 downto 0);
    signal IMA116_3638 : std_logic_vector(7 downto 0);
    signal IMA117_3648 : std_logic_vector(7 downto 0);
    signal IMA118_3658 : std_logic_vector(7 downto 0);
    signal IMA119_3668 : std_logic_vector(7 downto 0);
    signal IMA11_2588 : std_logic_vector(7 downto 0);
    signal IMA120_3678 : std_logic_vector(7 downto 0);
    signal IMA121_3688 : std_logic_vector(7 downto 0);
    signal IMA122_3698 : std_logic_vector(7 downto 0);
    signal IMA123_3708 : std_logic_vector(7 downto 0);
    signal IMA124_3718 : std_logic_vector(7 downto 0);
    signal IMA125_3728 : std_logic_vector(7 downto 0);
    signal IMA126_3738 : std_logic_vector(7 downto 0);
    signal IMA127_3748 : std_logic_vector(7 downto 0);
    signal IMA12_2598 : std_logic_vector(7 downto 0);
    signal IMA13_2608 : std_logic_vector(7 downto 0);
    signal IMA14_2618 : std_logic_vector(7 downto 0);
    signal IMA15_2628 : std_logic_vector(7 downto 0);
    signal IMA16_2638 : std_logic_vector(7 downto 0);
    signal IMA17_2648 : std_logic_vector(7 downto 0);
    signal IMA18_2658 : std_logic_vector(7 downto 0);
    signal IMA19_2668 : std_logic_vector(7 downto 0);
    signal IMA1_2488 : std_logic_vector(7 downto 0);
    signal IMA20_2678 : std_logic_vector(7 downto 0);
    signal IMA21_2688 : std_logic_vector(7 downto 0);
    signal IMA22_2698 : std_logic_vector(7 downto 0);
    signal IMA23_2708 : std_logic_vector(7 downto 0);
    signal IMA24_2718 : std_logic_vector(7 downto 0);
    signal IMA25_2728 : std_logic_vector(7 downto 0);
    signal IMA26_2738 : std_logic_vector(7 downto 0);
    signal IMA27_2748 : std_logic_vector(7 downto 0);
    signal IMA28_2758 : std_logic_vector(7 downto 0);
    signal IMA29_2768 : std_logic_vector(7 downto 0);
    signal IMA2_2498 : std_logic_vector(7 downto 0);
    signal IMA30_2778 : std_logic_vector(7 downto 0);
    signal IMA31_2788 : std_logic_vector(7 downto 0);
    signal IMA32_2798 : std_logic_vector(7 downto 0);
    signal IMA33_2808 : std_logic_vector(7 downto 0);
    signal IMA34_2818 : std_logic_vector(7 downto 0);
    signal IMA35_2828 : std_logic_vector(7 downto 0);
    signal IMA36_2838 : std_logic_vector(7 downto 0);
    signal IMA37_2848 : std_logic_vector(7 downto 0);
    signal IMA38_2858 : std_logic_vector(7 downto 0);
    signal IMA39_2868 : std_logic_vector(7 downto 0);
    signal IMA3_2508 : std_logic_vector(7 downto 0);
    signal IMA40_2878 : std_logic_vector(7 downto 0);
    signal IMA41_2888 : std_logic_vector(7 downto 0);
    signal IMA42_2898 : std_logic_vector(7 downto 0);
    signal IMA43_2908 : std_logic_vector(7 downto 0);
    signal IMA44_2918 : std_logic_vector(7 downto 0);
    signal IMA45_2928 : std_logic_vector(7 downto 0);
    signal IMA46_2938 : std_logic_vector(7 downto 0);
    signal IMA47_2948 : std_logic_vector(7 downto 0);
    signal IMA48_2958 : std_logic_vector(7 downto 0);
    signal IMA49_2968 : std_logic_vector(7 downto 0);
    signal IMA4_2518 : std_logic_vector(7 downto 0);
    signal IMA50_2978 : std_logic_vector(7 downto 0);
    signal IMA51_2988 : std_logic_vector(7 downto 0);
    signal IMA52_2998 : std_logic_vector(7 downto 0);
    signal IMA53_3008 : std_logic_vector(7 downto 0);
    signal IMA54_3018 : std_logic_vector(7 downto 0);
    signal IMA55_3028 : std_logic_vector(7 downto 0);
    signal IMA56_3038 : std_logic_vector(7 downto 0);
    signal IMA57_3048 : std_logic_vector(7 downto 0);
    signal IMA58_3058 : std_logic_vector(7 downto 0);
    signal IMA59_3068 : std_logic_vector(7 downto 0);
    signal IMA5_2528 : std_logic_vector(7 downto 0);
    signal IMA60_3078 : std_logic_vector(7 downto 0);
    signal IMA61_3088 : std_logic_vector(7 downto 0);
    signal IMA62_3098 : std_logic_vector(7 downto 0);
    signal IMA63_3108 : std_logic_vector(7 downto 0);
    signal IMA64_3118 : std_logic_vector(7 downto 0);
    signal IMA65_3128 : std_logic_vector(7 downto 0);
    signal IMA66_3138 : std_logic_vector(7 downto 0);
    signal IMA67_3148 : std_logic_vector(7 downto 0);
    signal IMA68_3158 : std_logic_vector(7 downto 0);
    signal IMA69_3168 : std_logic_vector(7 downto 0);
    signal IMA6_2538 : std_logic_vector(7 downto 0);
    signal IMA70_3178 : std_logic_vector(7 downto 0);
    signal IMA71_3188 : std_logic_vector(7 downto 0);
    signal IMA72_3198 : std_logic_vector(7 downto 0);
    signal IMA73_3208 : std_logic_vector(7 downto 0);
    signal IMA74_3218 : std_logic_vector(7 downto 0);
    signal IMA75_3228 : std_logic_vector(7 downto 0);
    signal IMA76_3238 : std_logic_vector(7 downto 0);
    signal IMA77_3248 : std_logic_vector(7 downto 0);
    signal IMA78_3258 : std_logic_vector(7 downto 0);
    signal IMA79_3268 : std_logic_vector(7 downto 0);
    signal IMA7_2548 : std_logic_vector(7 downto 0);
    signal IMA80_3278 : std_logic_vector(7 downto 0);
    signal IMA81_3288 : std_logic_vector(7 downto 0);
    signal IMA82_3298 : std_logic_vector(7 downto 0);
    signal IMA83_3308 : std_logic_vector(7 downto 0);
    signal IMA84_3318 : std_logic_vector(7 downto 0);
    signal IMA85_3328 : std_logic_vector(7 downto 0);
    signal IMA86_3338 : std_logic_vector(7 downto 0);
    signal IMA87_3348 : std_logic_vector(7 downto 0);
    signal IMA88_3358 : std_logic_vector(7 downto 0);
    signal IMA89_3368 : std_logic_vector(7 downto 0);
    signal IMA8_2558 : std_logic_vector(7 downto 0);
    signal IMA90_3378 : std_logic_vector(7 downto 0);
    signal IMA91_3388 : std_logic_vector(7 downto 0);
    signal IMA92_3398 : std_logic_vector(7 downto 0);
    signal IMA93_3408 : std_logic_vector(7 downto 0);
    signal IMA94_3418 : std_logic_vector(7 downto 0);
    signal IMA95_3428 : std_logic_vector(7 downto 0);
    signal IMA96_3438 : std_logic_vector(7 downto 0);
    signal IMA97_3448 : std_logic_vector(7 downto 0);
    signal IMA98_3458 : std_logic_vector(7 downto 0);
    signal IMA99_3468 : std_logic_vector(7 downto 0);
    signal IMA9_2568 : std_logic_vector(7 downto 0);
    signal IMB0_3756 : std_logic_vector(7 downto 0);
    signal IMB10_3836 : std_logic_vector(7 downto 0);
    signal IMB11_3844 : std_logic_vector(7 downto 0);
    signal IMB12_3852 : std_logic_vector(7 downto 0);
    signal IMB13_3860 : std_logic_vector(7 downto 0);
    signal IMB14_3868 : std_logic_vector(7 downto 0);
    signal IMB15_3876 : std_logic_vector(7 downto 0);
    signal IMB16_3884 : std_logic_vector(7 downto 0);
    signal IMB17_3892 : std_logic_vector(7 downto 0);
    signal IMB18_3900 : std_logic_vector(7 downto 0);
    signal IMB19_3908 : std_logic_vector(7 downto 0);
    signal IMB1_3764 : std_logic_vector(7 downto 0);
    signal IMB20_3916 : std_logic_vector(7 downto 0);
    signal IMB21_3924 : std_logic_vector(7 downto 0);
    signal IMB22_3932 : std_logic_vector(7 downto 0);
    signal IMB23_3940 : std_logic_vector(7 downto 0);
    signal IMB24_3948 : std_logic_vector(7 downto 0);
    signal IMB25_3956 : std_logic_vector(7 downto 0);
    signal IMB26_3964 : std_logic_vector(7 downto 0);
    signal IMB27_3972 : std_logic_vector(7 downto 0);
    signal IMB28_3980 : std_logic_vector(7 downto 0);
    signal IMB29_3988 : std_logic_vector(7 downto 0);
    signal IMB2_3772 : std_logic_vector(7 downto 0);
    signal IMB30_3996 : std_logic_vector(7 downto 0);
    signal IMB31_4004 : std_logic_vector(7 downto 0);
    signal IMB32_4012 : std_logic_vector(7 downto 0);
    signal IMB33_4020 : std_logic_vector(7 downto 0);
    signal IMB34_4028 : std_logic_vector(7 downto 0);
    signal IMB35_4036 : std_logic_vector(7 downto 0);
    signal IMB36_4044 : std_logic_vector(7 downto 0);
    signal IMB37_4052 : std_logic_vector(7 downto 0);
    signal IMB38_4060 : std_logic_vector(7 downto 0);
    signal IMB39_4068 : std_logic_vector(7 downto 0);
    signal IMB3_3780 : std_logic_vector(7 downto 0);
    signal IMB40_4076 : std_logic_vector(7 downto 0);
    signal IMB41_4084 : std_logic_vector(7 downto 0);
    signal IMB42_4092 : std_logic_vector(7 downto 0);
    signal IMB43_4100 : std_logic_vector(7 downto 0);
    signal IMB44_4108 : std_logic_vector(7 downto 0);
    signal IMB45_4116 : std_logic_vector(7 downto 0);
    signal IMB46_4124 : std_logic_vector(7 downto 0);
    signal IMB47_4132 : std_logic_vector(7 downto 0);
    signal IMB48_4140 : std_logic_vector(7 downto 0);
    signal IMB49_4148 : std_logic_vector(7 downto 0);
    signal IMB4_3788 : std_logic_vector(7 downto 0);
    signal IMB50_4156 : std_logic_vector(7 downto 0);
    signal IMB51_4164 : std_logic_vector(7 downto 0);
    signal IMB52_4172 : std_logic_vector(7 downto 0);
    signal IMB53_4180 : std_logic_vector(7 downto 0);
    signal IMB54_4188 : std_logic_vector(7 downto 0);
    signal IMB55_4196 : std_logic_vector(7 downto 0);
    signal IMB56_4204 : std_logic_vector(7 downto 0);
    signal IMB57_4212 : std_logic_vector(7 downto 0);
    signal IMB58_4220 : std_logic_vector(7 downto 0);
    signal IMB59_4228 : std_logic_vector(7 downto 0);
    signal IMB5_3796 : std_logic_vector(7 downto 0);
    signal IMB60_4236 : std_logic_vector(7 downto 0);
    signal IMB61_4244 : std_logic_vector(7 downto 0);
    signal IMB62_4252 : std_logic_vector(7 downto 0);
    signal IMB63_4260 : std_logic_vector(7 downto 0);
    signal IMB6_3804 : std_logic_vector(7 downto 0);
    signal IMB7_3812 : std_logic_vector(7 downto 0);
    signal IMB8_3820 : std_logic_vector(7 downto 0);
    signal IMB9_3828 : std_logic_vector(7 downto 0);
    signal IMC0_4268 : std_logic_vector(7 downto 0);
    signal IMC10_4348 : std_logic_vector(7 downto 0);
    signal IMC11_4356 : std_logic_vector(7 downto 0);
    signal IMC12_4364 : std_logic_vector(7 downto 0);
    signal IMC13_4372 : std_logic_vector(7 downto 0);
    signal IMC14_4380 : std_logic_vector(7 downto 0);
    signal IMC15_4388 : std_logic_vector(7 downto 0);
    signal IMC16_4396 : std_logic_vector(7 downto 0);
    signal IMC17_4404 : std_logic_vector(7 downto 0);
    signal IMC18_4412 : std_logic_vector(7 downto 0);
    signal IMC19_4420 : std_logic_vector(7 downto 0);
    signal IMC1_4276 : std_logic_vector(7 downto 0);
    signal IMC20_4428 : std_logic_vector(7 downto 0);
    signal IMC21_4436 : std_logic_vector(7 downto 0);
    signal IMC22_4444 : std_logic_vector(7 downto 0);
    signal IMC23_4452 : std_logic_vector(7 downto 0);
    signal IMC24_4460 : std_logic_vector(7 downto 0);
    signal IMC25_4468 : std_logic_vector(7 downto 0);
    signal IMC26_4476 : std_logic_vector(7 downto 0);
    signal IMC27_4484 : std_logic_vector(7 downto 0);
    signal IMC28_4492 : std_logic_vector(7 downto 0);
    signal IMC29_4500 : std_logic_vector(7 downto 0);
    signal IMC2_4284 : std_logic_vector(7 downto 0);
    signal IMC30_4508 : std_logic_vector(7 downto 0);
    signal IMC31_4516 : std_logic_vector(7 downto 0);
    signal IMC3_4292 : std_logic_vector(7 downto 0);
    signal IMC4_4300 : std_logic_vector(7 downto 0);
    signal IMC5_4308 : std_logic_vector(7 downto 0);
    signal IMC6_4316 : std_logic_vector(7 downto 0);
    signal IMC7_4324 : std_logic_vector(7 downto 0);
    signal IMC8_4332 : std_logic_vector(7 downto 0);
    signal IMC9_4340 : std_logic_vector(7 downto 0);
    signal IMD0_4524 : std_logic_vector(7 downto 0);
    signal IMD10_4604 : std_logic_vector(7 downto 0);
    signal IMD11_4612 : std_logic_vector(7 downto 0);
    signal IMD12_4620 : std_logic_vector(7 downto 0);
    signal IMD13_4628 : std_logic_vector(7 downto 0);
    signal IMD14_4636 : std_logic_vector(7 downto 0);
    signal IMD15_4644 : std_logic_vector(7 downto 0);
    signal IMD1_4532 : std_logic_vector(7 downto 0);
    signal IMD2_4540 : std_logic_vector(7 downto 0);
    signal IMD3_4548 : std_logic_vector(7 downto 0);
    signal IMD4_4556 : std_logic_vector(7 downto 0);
    signal IMD5_4564 : std_logic_vector(7 downto 0);
    signal IMD6_4572 : std_logic_vector(7 downto 0);
    signal IMD7_4580 : std_logic_vector(7 downto 0);
    signal IMD8_4588 : std_logic_vector(7 downto 0);
    signal IMD9_4596 : std_logic_vector(7 downto 0);
    signal IME0_4652 : std_logic_vector(7 downto 0);
    signal IME1_4660 : std_logic_vector(7 downto 0);
    signal IME2_4668 : std_logic_vector(7 downto 0);
    signal IME3_4676 : std_logic_vector(7 downto 0);
    signal IME4_4684 : std_logic_vector(7 downto 0);
    signal IME5_4692 : std_logic_vector(7 downto 0);
    signal IME6_4700 : std_logic_vector(7 downto 0);
    signal IME7_4708 : std_logic_vector(7 downto 0);
    signal IMF0_4716 : std_logic_vector(7 downto 0);
    signal IMF1_4724 : std_logic_vector(7 downto 0);
    signal IMF2_4732 : std_logic_vector(7 downto 0);
    signal IMF3_4740 : std_logic_vector(7 downto 0);
    signal IMG0_4748 : std_logic_vector(7 downto 0);
    signal IMG1_4756 : std_logic_vector(7 downto 0);
    signal konst_2471_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2481_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2491_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2501_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2511_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2521_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2531_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2541_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2551_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2561_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2571_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2581_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2591_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2601_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2611_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2621_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2631_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2641_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2651_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2661_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2671_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2681_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2691_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2701_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2711_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2721_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2731_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2741_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2751_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2761_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2771_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2781_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2791_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2801_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2811_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2821_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2831_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2841_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2851_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2861_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2871_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2881_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2891_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2901_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2911_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2921_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2931_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2941_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2951_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2961_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2971_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2981_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2991_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3001_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3011_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3021_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3031_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3041_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3051_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3061_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3071_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3081_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3091_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3101_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3111_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3121_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3131_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3141_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3151_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3161_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3171_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3181_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3191_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3201_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3211_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3221_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3231_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3241_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3251_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3261_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3271_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3281_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3291_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3301_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3311_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3321_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3331_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3341_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3351_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3361_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3371_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3381_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3391_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3401_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3411_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3421_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3431_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3441_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3451_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3461_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3471_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3481_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3491_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3501_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3511_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3521_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3531_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3541_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3551_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3561_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3571_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3581_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3591_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3601_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3611_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3621_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3631_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3641_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3651_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3661_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3671_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3681_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3691_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3701_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3711_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3721_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3731_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3741_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3751_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3759_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3767_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3775_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3783_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3791_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3799_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3807_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3815_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3823_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3831_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3839_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3847_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3855_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3863_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3871_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3879_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3887_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3895_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3903_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3911_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3919_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3927_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3935_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3943_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3951_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3959_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3967_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3975_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3983_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3991_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3999_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4007_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4015_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4023_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4031_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4039_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4047_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4055_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4063_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4071_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4079_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4087_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4095_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4103_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4111_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4119_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4127_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4135_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4143_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4151_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4159_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4167_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4175_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4183_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4191_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4199_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4207_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4215_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4223_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4231_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4239_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4247_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4255_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4263_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4271_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4279_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4287_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4295_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4303_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4311_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4319_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4327_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4335_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4343_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4351_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4359_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4367_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4375_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4383_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4391_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4399_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4407_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4415_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4423_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4431_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4439_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4447_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4455_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4463_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4471_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4479_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4487_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4495_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4503_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4511_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4519_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4527_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4535_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4543_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4551_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4559_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4567_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4575_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4583_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4591_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4599_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4607_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4615_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4623_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4631_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4639_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4647_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4655_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4663_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4671_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4679_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4687_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4695_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4703_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4711_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4719_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4727_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4735_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4743_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4751_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4759_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2474_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2476_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2484_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2486_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2494_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2496_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2504_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2506_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2514_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2516_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2524_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2526_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2534_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2536_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2544_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2546_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2554_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2556_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2564_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2566_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2574_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2576_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2584_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2586_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2594_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2596_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2604_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2606_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2614_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2616_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2624_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2626_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2634_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2636_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2644_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2646_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2654_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2656_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2664_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2666_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2674_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2676_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2684_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2686_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2694_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2696_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2704_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2706_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2714_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2716_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2724_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2726_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2734_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2736_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2744_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2746_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2754_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2756_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2764_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2766_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2774_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2776_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2784_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2786_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2794_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2796_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2804_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2806_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2814_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2816_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2824_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2826_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2834_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2836_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2844_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2846_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2854_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2856_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2864_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2866_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2874_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2876_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2884_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2886_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2894_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2896_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2904_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2906_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2914_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2916_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2924_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2926_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2934_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2936_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2944_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2946_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2954_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2956_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2964_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2966_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2974_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2976_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2984_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2986_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2994_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2996_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3004_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3006_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3014_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3016_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3024_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3026_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3034_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3036_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3044_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3046_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3054_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3056_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3064_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3066_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3074_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3076_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3084_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3086_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3094_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3096_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3104_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3106_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3114_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3116_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3124_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3126_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3134_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3136_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3144_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3146_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3154_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3156_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3164_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3166_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3174_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3176_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3184_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3186_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3194_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3196_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3204_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3206_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3214_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3216_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3224_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3226_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3234_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3236_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3244_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3246_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3254_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3256_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3264_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3266_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3274_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3276_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3284_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3286_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3294_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3296_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3304_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3306_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3314_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3316_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3324_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3326_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3334_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3336_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3344_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3346_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3354_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3356_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3364_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3366_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3374_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3376_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3384_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3386_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3394_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3396_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3404_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3406_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3414_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3416_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3424_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3426_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3434_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3436_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3444_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3446_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3454_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3456_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3464_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3466_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3474_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3476_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3484_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3486_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3494_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3496_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3504_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3506_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3514_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3516_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3524_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3526_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3534_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3536_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3544_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3546_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3554_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3556_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3564_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3566_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3574_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3576_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3584_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3586_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3594_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3596_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3604_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3606_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3614_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3616_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3624_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3626_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3634_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3636_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3644_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3646_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3654_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3656_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3664_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3666_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3674_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3676_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3684_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3686_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3694_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3696_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3704_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3706_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3714_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3716_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3724_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3726_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3734_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3736_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3744_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3746_wire_constant : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    konst_2471_wire_constant <= "00000000";
    konst_2481_wire_constant <= "00000000";
    konst_2491_wire_constant <= "00000000";
    konst_2501_wire_constant <= "00000000";
    konst_2511_wire_constant <= "00000000";
    konst_2521_wire_constant <= "00000000";
    konst_2531_wire_constant <= "00000000";
    konst_2541_wire_constant <= "00000000";
    konst_2551_wire_constant <= "00000000";
    konst_2561_wire_constant <= "00000000";
    konst_2571_wire_constant <= "00000000";
    konst_2581_wire_constant <= "00000000";
    konst_2591_wire_constant <= "00000000";
    konst_2601_wire_constant <= "00000000";
    konst_2611_wire_constant <= "00000000";
    konst_2621_wire_constant <= "00000000";
    konst_2631_wire_constant <= "00000000";
    konst_2641_wire_constant <= "00000000";
    konst_2651_wire_constant <= "00000000";
    konst_2661_wire_constant <= "00000000";
    konst_2671_wire_constant <= "00000000";
    konst_2681_wire_constant <= "00000000";
    konst_2691_wire_constant <= "00000000";
    konst_2701_wire_constant <= "00000000";
    konst_2711_wire_constant <= "00000000";
    konst_2721_wire_constant <= "00000000";
    konst_2731_wire_constant <= "00000000";
    konst_2741_wire_constant <= "00000000";
    konst_2751_wire_constant <= "00000000";
    konst_2761_wire_constant <= "00000000";
    konst_2771_wire_constant <= "00000000";
    konst_2781_wire_constant <= "00000000";
    konst_2791_wire_constant <= "00000000";
    konst_2801_wire_constant <= "00000000";
    konst_2811_wire_constant <= "00000000";
    konst_2821_wire_constant <= "00000000";
    konst_2831_wire_constant <= "00000000";
    konst_2841_wire_constant <= "00000000";
    konst_2851_wire_constant <= "00000000";
    konst_2861_wire_constant <= "00000000";
    konst_2871_wire_constant <= "00000000";
    konst_2881_wire_constant <= "00000000";
    konst_2891_wire_constant <= "00000000";
    konst_2901_wire_constant <= "00000000";
    konst_2911_wire_constant <= "00000000";
    konst_2921_wire_constant <= "00000000";
    konst_2931_wire_constant <= "00000000";
    konst_2941_wire_constant <= "00000000";
    konst_2951_wire_constant <= "00000000";
    konst_2961_wire_constant <= "00000000";
    konst_2971_wire_constant <= "00000000";
    konst_2981_wire_constant <= "00000000";
    konst_2991_wire_constant <= "00000000";
    konst_3001_wire_constant <= "00000000";
    konst_3011_wire_constant <= "00000000";
    konst_3021_wire_constant <= "00000000";
    konst_3031_wire_constant <= "00000000";
    konst_3041_wire_constant <= "00000000";
    konst_3051_wire_constant <= "00000000";
    konst_3061_wire_constant <= "00000000";
    konst_3071_wire_constant <= "00000000";
    konst_3081_wire_constant <= "00000000";
    konst_3091_wire_constant <= "00000000";
    konst_3101_wire_constant <= "00000000";
    konst_3111_wire_constant <= "00000000";
    konst_3121_wire_constant <= "00000000";
    konst_3131_wire_constant <= "00000000";
    konst_3141_wire_constant <= "00000000";
    konst_3151_wire_constant <= "00000000";
    konst_3161_wire_constant <= "00000000";
    konst_3171_wire_constant <= "00000000";
    konst_3181_wire_constant <= "00000000";
    konst_3191_wire_constant <= "00000000";
    konst_3201_wire_constant <= "00000000";
    konst_3211_wire_constant <= "00000000";
    konst_3221_wire_constant <= "00000000";
    konst_3231_wire_constant <= "00000000";
    konst_3241_wire_constant <= "00000000";
    konst_3251_wire_constant <= "00000000";
    konst_3261_wire_constant <= "00000000";
    konst_3271_wire_constant <= "00000000";
    konst_3281_wire_constant <= "00000000";
    konst_3291_wire_constant <= "00000000";
    konst_3301_wire_constant <= "00000000";
    konst_3311_wire_constant <= "00000000";
    konst_3321_wire_constant <= "00000000";
    konst_3331_wire_constant <= "00000000";
    konst_3341_wire_constant <= "00000000";
    konst_3351_wire_constant <= "00000000";
    konst_3361_wire_constant <= "00000000";
    konst_3371_wire_constant <= "00000000";
    konst_3381_wire_constant <= "00000000";
    konst_3391_wire_constant <= "00000000";
    konst_3401_wire_constant <= "00000000";
    konst_3411_wire_constant <= "00000000";
    konst_3421_wire_constant <= "00000000";
    konst_3431_wire_constant <= "00000000";
    konst_3441_wire_constant <= "00000000";
    konst_3451_wire_constant <= "00000000";
    konst_3461_wire_constant <= "00000000";
    konst_3471_wire_constant <= "00000000";
    konst_3481_wire_constant <= "00000000";
    konst_3491_wire_constant <= "00000000";
    konst_3501_wire_constant <= "00000000";
    konst_3511_wire_constant <= "00000000";
    konst_3521_wire_constant <= "00000000";
    konst_3531_wire_constant <= "00000000";
    konst_3541_wire_constant <= "00000000";
    konst_3551_wire_constant <= "00000000";
    konst_3561_wire_constant <= "00000000";
    konst_3571_wire_constant <= "00000000";
    konst_3581_wire_constant <= "00000000";
    konst_3591_wire_constant <= "00000000";
    konst_3601_wire_constant <= "00000000";
    konst_3611_wire_constant <= "00000000";
    konst_3621_wire_constant <= "00000000";
    konst_3631_wire_constant <= "00000000";
    konst_3641_wire_constant <= "00000000";
    konst_3651_wire_constant <= "00000000";
    konst_3661_wire_constant <= "00000000";
    konst_3671_wire_constant <= "00000000";
    konst_3681_wire_constant <= "00000000";
    konst_3691_wire_constant <= "00000000";
    konst_3701_wire_constant <= "00000000";
    konst_3711_wire_constant <= "00000000";
    konst_3721_wire_constant <= "00000000";
    konst_3731_wire_constant <= "00000000";
    konst_3741_wire_constant <= "00000000";
    konst_3751_wire_constant <= "00000001";
    konst_3759_wire_constant <= "00000001";
    konst_3767_wire_constant <= "00000001";
    konst_3775_wire_constant <= "00000001";
    konst_3783_wire_constant <= "00000001";
    konst_3791_wire_constant <= "00000001";
    konst_3799_wire_constant <= "00000001";
    konst_3807_wire_constant <= "00000001";
    konst_3815_wire_constant <= "00000001";
    konst_3823_wire_constant <= "00000001";
    konst_3831_wire_constant <= "00000001";
    konst_3839_wire_constant <= "00000001";
    konst_3847_wire_constant <= "00000001";
    konst_3855_wire_constant <= "00000001";
    konst_3863_wire_constant <= "00000001";
    konst_3871_wire_constant <= "00000001";
    konst_3879_wire_constant <= "00000001";
    konst_3887_wire_constant <= "00000001";
    konst_3895_wire_constant <= "00000001";
    konst_3903_wire_constant <= "00000001";
    konst_3911_wire_constant <= "00000001";
    konst_3919_wire_constant <= "00000001";
    konst_3927_wire_constant <= "00000001";
    konst_3935_wire_constant <= "00000001";
    konst_3943_wire_constant <= "00000001";
    konst_3951_wire_constant <= "00000001";
    konst_3959_wire_constant <= "00000001";
    konst_3967_wire_constant <= "00000001";
    konst_3975_wire_constant <= "00000001";
    konst_3983_wire_constant <= "00000001";
    konst_3991_wire_constant <= "00000001";
    konst_3999_wire_constant <= "00000001";
    konst_4007_wire_constant <= "00000001";
    konst_4015_wire_constant <= "00000001";
    konst_4023_wire_constant <= "00000001";
    konst_4031_wire_constant <= "00000001";
    konst_4039_wire_constant <= "00000001";
    konst_4047_wire_constant <= "00000001";
    konst_4055_wire_constant <= "00000001";
    konst_4063_wire_constant <= "00000001";
    konst_4071_wire_constant <= "00000001";
    konst_4079_wire_constant <= "00000001";
    konst_4087_wire_constant <= "00000001";
    konst_4095_wire_constant <= "00000001";
    konst_4103_wire_constant <= "00000001";
    konst_4111_wire_constant <= "00000001";
    konst_4119_wire_constant <= "00000001";
    konst_4127_wire_constant <= "00000001";
    konst_4135_wire_constant <= "00000001";
    konst_4143_wire_constant <= "00000001";
    konst_4151_wire_constant <= "00000001";
    konst_4159_wire_constant <= "00000001";
    konst_4167_wire_constant <= "00000001";
    konst_4175_wire_constant <= "00000001";
    konst_4183_wire_constant <= "00000001";
    konst_4191_wire_constant <= "00000001";
    konst_4199_wire_constant <= "00000001";
    konst_4207_wire_constant <= "00000001";
    konst_4215_wire_constant <= "00000001";
    konst_4223_wire_constant <= "00000001";
    konst_4231_wire_constant <= "00000001";
    konst_4239_wire_constant <= "00000001";
    konst_4247_wire_constant <= "00000001";
    konst_4255_wire_constant <= "00000001";
    konst_4263_wire_constant <= "00000010";
    konst_4271_wire_constant <= "00000010";
    konst_4279_wire_constant <= "00000010";
    konst_4287_wire_constant <= "00000010";
    konst_4295_wire_constant <= "00000010";
    konst_4303_wire_constant <= "00000010";
    konst_4311_wire_constant <= "00000010";
    konst_4319_wire_constant <= "00000010";
    konst_4327_wire_constant <= "00000010";
    konst_4335_wire_constant <= "00000010";
    konst_4343_wire_constant <= "00000010";
    konst_4351_wire_constant <= "00000010";
    konst_4359_wire_constant <= "00000010";
    konst_4367_wire_constant <= "00000010";
    konst_4375_wire_constant <= "00000010";
    konst_4383_wire_constant <= "00000010";
    konst_4391_wire_constant <= "00000010";
    konst_4399_wire_constant <= "00000010";
    konst_4407_wire_constant <= "00000010";
    konst_4415_wire_constant <= "00000010";
    konst_4423_wire_constant <= "00000010";
    konst_4431_wire_constant <= "00000010";
    konst_4439_wire_constant <= "00000010";
    konst_4447_wire_constant <= "00000010";
    konst_4455_wire_constant <= "00000010";
    konst_4463_wire_constant <= "00000010";
    konst_4471_wire_constant <= "00000010";
    konst_4479_wire_constant <= "00000010";
    konst_4487_wire_constant <= "00000010";
    konst_4495_wire_constant <= "00000010";
    konst_4503_wire_constant <= "00000010";
    konst_4511_wire_constant <= "00000010";
    konst_4519_wire_constant <= "00000011";
    konst_4527_wire_constant <= "00000011";
    konst_4535_wire_constant <= "00000011";
    konst_4543_wire_constant <= "00000011";
    konst_4551_wire_constant <= "00000011";
    konst_4559_wire_constant <= "00000011";
    konst_4567_wire_constant <= "00000011";
    konst_4575_wire_constant <= "00000011";
    konst_4583_wire_constant <= "00000011";
    konst_4591_wire_constant <= "00000011";
    konst_4599_wire_constant <= "00000011";
    konst_4607_wire_constant <= "00000011";
    konst_4615_wire_constant <= "00000011";
    konst_4623_wire_constant <= "00000011";
    konst_4631_wire_constant <= "00000011";
    konst_4639_wire_constant <= "00000011";
    konst_4647_wire_constant <= "00000100";
    konst_4655_wire_constant <= "00000100";
    konst_4663_wire_constant <= "00000100";
    konst_4671_wire_constant <= "00000100";
    konst_4679_wire_constant <= "00000100";
    konst_4687_wire_constant <= "00000100";
    konst_4695_wire_constant <= "00000100";
    konst_4703_wire_constant <= "00000100";
    konst_4711_wire_constant <= "00000101";
    konst_4719_wire_constant <= "00000101";
    konst_4727_wire_constant <= "00000101";
    konst_4735_wire_constant <= "00000101";
    konst_4743_wire_constant <= "00000110";
    konst_4751_wire_constant <= "00000110";
    konst_4759_wire_constant <= "00000111";
    type_cast_2474_wire_constant <= "00001001";
    type_cast_2476_wire_constant <= "01010010";
    type_cast_2484_wire_constant <= "11010101";
    type_cast_2486_wire_constant <= "01101010";
    type_cast_2494_wire_constant <= "00110110";
    type_cast_2496_wire_constant <= "00110000";
    type_cast_2504_wire_constant <= "00111000";
    type_cast_2506_wire_constant <= "10100101";
    type_cast_2514_wire_constant <= "01000000";
    type_cast_2516_wire_constant <= "10111111";
    type_cast_2524_wire_constant <= "10011110";
    type_cast_2526_wire_constant <= "10100011";
    type_cast_2534_wire_constant <= "11110011";
    type_cast_2536_wire_constant <= "10000001";
    type_cast_2544_wire_constant <= "11111011";
    type_cast_2546_wire_constant <= "11010111";
    type_cast_2554_wire_constant <= "11100011";
    type_cast_2556_wire_constant <= "01111100";
    type_cast_2564_wire_constant <= "10000010";
    type_cast_2566_wire_constant <= "00111001";
    type_cast_2574_wire_constant <= "00101111";
    type_cast_2576_wire_constant <= "10011011";
    type_cast_2584_wire_constant <= "10000111";
    type_cast_2586_wire_constant <= "11111111";
    type_cast_2594_wire_constant <= "10001110";
    type_cast_2596_wire_constant <= "00110100";
    type_cast_2604_wire_constant <= "01000100";
    type_cast_2606_wire_constant <= "01000011";
    type_cast_2614_wire_constant <= "11011110";
    type_cast_2616_wire_constant <= "11000100";
    type_cast_2624_wire_constant <= "11001011";
    type_cast_2626_wire_constant <= "11101001";
    type_cast_2634_wire_constant <= "01111011";
    type_cast_2636_wire_constant <= "01010100";
    type_cast_2644_wire_constant <= "00110010";
    type_cast_2646_wire_constant <= "10010100";
    type_cast_2654_wire_constant <= "11000010";
    type_cast_2656_wire_constant <= "10100110";
    type_cast_2664_wire_constant <= "00111101";
    type_cast_2666_wire_constant <= "00100011";
    type_cast_2674_wire_constant <= "01001100";
    type_cast_2676_wire_constant <= "11101110";
    type_cast_2684_wire_constant <= "00001011";
    type_cast_2686_wire_constant <= "10010101";
    type_cast_2694_wire_constant <= "11111010";
    type_cast_2696_wire_constant <= "01000010";
    type_cast_2704_wire_constant <= "01001110";
    type_cast_2706_wire_constant <= "11000011";
    type_cast_2714_wire_constant <= "00101110";
    type_cast_2716_wire_constant <= "00001000";
    type_cast_2724_wire_constant <= "01100110";
    type_cast_2726_wire_constant <= "10100001";
    type_cast_2734_wire_constant <= "11011001";
    type_cast_2736_wire_constant <= "00101000";
    type_cast_2744_wire_constant <= "10110010";
    type_cast_2746_wire_constant <= "00100100";
    type_cast_2754_wire_constant <= "01011011";
    type_cast_2756_wire_constant <= "01110110";
    type_cast_2764_wire_constant <= "01001001";
    type_cast_2766_wire_constant <= "10100010";
    type_cast_2774_wire_constant <= "10001011";
    type_cast_2776_wire_constant <= "01101101";
    type_cast_2784_wire_constant <= "00100101";
    type_cast_2786_wire_constant <= "11010001";
    type_cast_2794_wire_constant <= "11111000";
    type_cast_2796_wire_constant <= "01110010";
    type_cast_2804_wire_constant <= "01100100";
    type_cast_2806_wire_constant <= "11110110";
    type_cast_2814_wire_constant <= "01101000";
    type_cast_2816_wire_constant <= "10000110";
    type_cast_2824_wire_constant <= "00010110";
    type_cast_2826_wire_constant <= "10011000";
    type_cast_2834_wire_constant <= "10100100";
    type_cast_2836_wire_constant <= "11010100";
    type_cast_2844_wire_constant <= "11001100";
    type_cast_2846_wire_constant <= "01011100";
    type_cast_2854_wire_constant <= "01100101";
    type_cast_2856_wire_constant <= "01011101";
    type_cast_2864_wire_constant <= "10010010";
    type_cast_2866_wire_constant <= "10110110";
    type_cast_2874_wire_constant <= "01110000";
    type_cast_2876_wire_constant <= "01101100";
    type_cast_2884_wire_constant <= "01010000";
    type_cast_2886_wire_constant <= "01001000";
    type_cast_2894_wire_constant <= "11101101";
    type_cast_2896_wire_constant <= "11111101";
    type_cast_2904_wire_constant <= "11011010";
    type_cast_2906_wire_constant <= "10111001";
    type_cast_2914_wire_constant <= "00010101";
    type_cast_2916_wire_constant <= "01011110";
    type_cast_2924_wire_constant <= "01010111";
    type_cast_2926_wire_constant <= "01000110";
    type_cast_2934_wire_constant <= "10001101";
    type_cast_2936_wire_constant <= "10100111";
    type_cast_2944_wire_constant <= "10000100";
    type_cast_2946_wire_constant <= "10011101";
    type_cast_2954_wire_constant <= "11011000";
    type_cast_2956_wire_constant <= "10010000";
    type_cast_2964_wire_constant <= "00000000";
    type_cast_2966_wire_constant <= "10101011";
    type_cast_2974_wire_constant <= "10111100";
    type_cast_2976_wire_constant <= "10001100";
    type_cast_2984_wire_constant <= "00001010";
    type_cast_2986_wire_constant <= "11010011";
    type_cast_2994_wire_constant <= "11100100";
    type_cast_2996_wire_constant <= "11110111";
    type_cast_3004_wire_constant <= "00000101";
    type_cast_3006_wire_constant <= "01011000";
    type_cast_3014_wire_constant <= "10110011";
    type_cast_3016_wire_constant <= "10111000";
    type_cast_3024_wire_constant <= "00000110";
    type_cast_3026_wire_constant <= "01000101";
    type_cast_3034_wire_constant <= "00101100";
    type_cast_3036_wire_constant <= "11010000";
    type_cast_3044_wire_constant <= "10001111";
    type_cast_3046_wire_constant <= "00011110";
    type_cast_3054_wire_constant <= "00111111";
    type_cast_3056_wire_constant <= "11001010";
    type_cast_3064_wire_constant <= "00000010";
    type_cast_3066_wire_constant <= "00001111";
    type_cast_3074_wire_constant <= "10101111";
    type_cast_3076_wire_constant <= "11000001";
    type_cast_3084_wire_constant <= "00000011";
    type_cast_3086_wire_constant <= "10111101";
    type_cast_3094_wire_constant <= "00010011";
    type_cast_3096_wire_constant <= "00000001";
    type_cast_3104_wire_constant <= "01101011";
    type_cast_3106_wire_constant <= "10001010";
    type_cast_3114_wire_constant <= "10010001";
    type_cast_3116_wire_constant <= "00111010";
    type_cast_3124_wire_constant <= "01000001";
    type_cast_3126_wire_constant <= "00010001";
    type_cast_3134_wire_constant <= "01100111";
    type_cast_3136_wire_constant <= "01001111";
    type_cast_3144_wire_constant <= "11101010";
    type_cast_3146_wire_constant <= "11011100";
    type_cast_3154_wire_constant <= "11110010";
    type_cast_3156_wire_constant <= "10010111";
    type_cast_3164_wire_constant <= "11001110";
    type_cast_3166_wire_constant <= "11001111";
    type_cast_3174_wire_constant <= "10110100";
    type_cast_3176_wire_constant <= "11110000";
    type_cast_3184_wire_constant <= "01110011";
    type_cast_3186_wire_constant <= "11100110";
    type_cast_3194_wire_constant <= "10101100";
    type_cast_3196_wire_constant <= "10010110";
    type_cast_3204_wire_constant <= "00100010";
    type_cast_3206_wire_constant <= "01110100";
    type_cast_3214_wire_constant <= "10101101";
    type_cast_3216_wire_constant <= "11100111";
    type_cast_3224_wire_constant <= "10000101";
    type_cast_3226_wire_constant <= "00110101";
    type_cast_3234_wire_constant <= "11111001";
    type_cast_3236_wire_constant <= "11100010";
    type_cast_3244_wire_constant <= "11101000";
    type_cast_3246_wire_constant <= "00110111";
    type_cast_3254_wire_constant <= "01110101";
    type_cast_3256_wire_constant <= "00011100";
    type_cast_3264_wire_constant <= "01101110";
    type_cast_3266_wire_constant <= "11011111";
    type_cast_3274_wire_constant <= "11110001";
    type_cast_3276_wire_constant <= "01000111";
    type_cast_3284_wire_constant <= "01110001";
    type_cast_3286_wire_constant <= "00011010";
    type_cast_3294_wire_constant <= "00101001";
    type_cast_3296_wire_constant <= "00011101";
    type_cast_3304_wire_constant <= "10001001";
    type_cast_3306_wire_constant <= "11000101";
    type_cast_3314_wire_constant <= "10110111";
    type_cast_3316_wire_constant <= "01101111";
    type_cast_3324_wire_constant <= "00001110";
    type_cast_3326_wire_constant <= "01100010";
    type_cast_3334_wire_constant <= "00011000";
    type_cast_3336_wire_constant <= "10101010";
    type_cast_3344_wire_constant <= "00011011";
    type_cast_3346_wire_constant <= "10111110";
    type_cast_3354_wire_constant <= "01010110";
    type_cast_3356_wire_constant <= "11111100";
    type_cast_3364_wire_constant <= "01001011";
    type_cast_3366_wire_constant <= "00111110";
    type_cast_3374_wire_constant <= "11010010";
    type_cast_3376_wire_constant <= "11000110";
    type_cast_3384_wire_constant <= "00100000";
    type_cast_3386_wire_constant <= "01111001";
    type_cast_3394_wire_constant <= "11011011";
    type_cast_3396_wire_constant <= "10011010";
    type_cast_3404_wire_constant <= "11111110";
    type_cast_3406_wire_constant <= "11000000";
    type_cast_3414_wire_constant <= "11001101";
    type_cast_3416_wire_constant <= "01111000";
    type_cast_3424_wire_constant <= "11110100";
    type_cast_3426_wire_constant <= "01011010";
    type_cast_3434_wire_constant <= "11011101";
    type_cast_3436_wire_constant <= "00011111";
    type_cast_3444_wire_constant <= "00110011";
    type_cast_3446_wire_constant <= "10101000";
    type_cast_3454_wire_constant <= "00000111";
    type_cast_3456_wire_constant <= "10001000";
    type_cast_3464_wire_constant <= "00110001";
    type_cast_3466_wire_constant <= "11000111";
    type_cast_3474_wire_constant <= "00010010";
    type_cast_3476_wire_constant <= "10110001";
    type_cast_3484_wire_constant <= "01011001";
    type_cast_3486_wire_constant <= "00010000";
    type_cast_3494_wire_constant <= "10000000";
    type_cast_3496_wire_constant <= "00100111";
    type_cast_3504_wire_constant <= "01011111";
    type_cast_3506_wire_constant <= "11101100";
    type_cast_3514_wire_constant <= "01010001";
    type_cast_3516_wire_constant <= "01100000";
    type_cast_3524_wire_constant <= "10101001";
    type_cast_3526_wire_constant <= "01111111";
    type_cast_3534_wire_constant <= "10110101";
    type_cast_3536_wire_constant <= "00011001";
    type_cast_3544_wire_constant <= "00001101";
    type_cast_3546_wire_constant <= "01001010";
    type_cast_3554_wire_constant <= "11100101";
    type_cast_3556_wire_constant <= "00101101";
    type_cast_3564_wire_constant <= "10011111";
    type_cast_3566_wire_constant <= "01111010";
    type_cast_3574_wire_constant <= "11001001";
    type_cast_3576_wire_constant <= "10010011";
    type_cast_3584_wire_constant <= "11101111";
    type_cast_3586_wire_constant <= "10011100";
    type_cast_3594_wire_constant <= "11100000";
    type_cast_3596_wire_constant <= "10100000";
    type_cast_3604_wire_constant <= "01001101";
    type_cast_3606_wire_constant <= "00111011";
    type_cast_3614_wire_constant <= "00101010";
    type_cast_3616_wire_constant <= "10101110";
    type_cast_3624_wire_constant <= "10110000";
    type_cast_3626_wire_constant <= "11110101";
    type_cast_3634_wire_constant <= "11101011";
    type_cast_3636_wire_constant <= "11001000";
    type_cast_3644_wire_constant <= "00111100";
    type_cast_3646_wire_constant <= "10111011";
    type_cast_3654_wire_constant <= "01010011";
    type_cast_3656_wire_constant <= "10000011";
    type_cast_3664_wire_constant <= "01100001";
    type_cast_3666_wire_constant <= "10011001";
    type_cast_3674_wire_constant <= "00101011";
    type_cast_3676_wire_constant <= "00010111";
    type_cast_3684_wire_constant <= "01111110";
    type_cast_3686_wire_constant <= "00000100";
    type_cast_3694_wire_constant <= "01110111";
    type_cast_3696_wire_constant <= "10111010";
    type_cast_3704_wire_constant <= "00100110";
    type_cast_3706_wire_constant <= "11010110";
    type_cast_3714_wire_constant <= "01101001";
    type_cast_3716_wire_constant <= "11100001";
    type_cast_3724_wire_constant <= "01100011";
    type_cast_3726_wire_constant <= "00010100";
    type_cast_3734_wire_constant <= "00100001";
    type_cast_3736_wire_constant <= "01010101";
    type_cast_3744_wire_constant <= "01111101";
    type_cast_3746_wire_constant <= "00001100";
    -- flow-through select operator MUX_2477_inst
    IMA0_2478 <= type_cast_2474_wire_constant when (BITSEL_u8_u1_2472_wire(0) /=  '0') else type_cast_2476_wire_constant;
    -- flow-through select operator MUX_2487_inst
    IMA1_2488 <= type_cast_2484_wire_constant when (BITSEL_u8_u1_2482_wire(0) /=  '0') else type_cast_2486_wire_constant;
    -- flow-through select operator MUX_2497_inst
    IMA2_2498 <= type_cast_2494_wire_constant when (BITSEL_u8_u1_2492_wire(0) /=  '0') else type_cast_2496_wire_constant;
    -- flow-through select operator MUX_2507_inst
    IMA3_2508 <= type_cast_2504_wire_constant when (BITSEL_u8_u1_2502_wire(0) /=  '0') else type_cast_2506_wire_constant;
    -- flow-through select operator MUX_2517_inst
    IMA4_2518 <= type_cast_2514_wire_constant when (BITSEL_u8_u1_2512_wire(0) /=  '0') else type_cast_2516_wire_constant;
    -- flow-through select operator MUX_2527_inst
    IMA5_2528 <= type_cast_2524_wire_constant when (BITSEL_u8_u1_2522_wire(0) /=  '0') else type_cast_2526_wire_constant;
    -- flow-through select operator MUX_2537_inst
    IMA6_2538 <= type_cast_2534_wire_constant when (BITSEL_u8_u1_2532_wire(0) /=  '0') else type_cast_2536_wire_constant;
    -- flow-through select operator MUX_2547_inst
    IMA7_2548 <= type_cast_2544_wire_constant when (BITSEL_u8_u1_2542_wire(0) /=  '0') else type_cast_2546_wire_constant;
    -- flow-through select operator MUX_2557_inst
    IMA8_2558 <= type_cast_2554_wire_constant when (BITSEL_u8_u1_2552_wire(0) /=  '0') else type_cast_2556_wire_constant;
    -- flow-through select operator MUX_2567_inst
    IMA9_2568 <= type_cast_2564_wire_constant when (BITSEL_u8_u1_2562_wire(0) /=  '0') else type_cast_2566_wire_constant;
    -- flow-through select operator MUX_2577_inst
    IMA10_2578 <= type_cast_2574_wire_constant when (BITSEL_u8_u1_2572_wire(0) /=  '0') else type_cast_2576_wire_constant;
    -- flow-through select operator MUX_2587_inst
    IMA11_2588 <= type_cast_2584_wire_constant when (BITSEL_u8_u1_2582_wire(0) /=  '0') else type_cast_2586_wire_constant;
    -- flow-through select operator MUX_2597_inst
    IMA12_2598 <= type_cast_2594_wire_constant when (BITSEL_u8_u1_2592_wire(0) /=  '0') else type_cast_2596_wire_constant;
    -- flow-through select operator MUX_2607_inst
    IMA13_2608 <= type_cast_2604_wire_constant when (BITSEL_u8_u1_2602_wire(0) /=  '0') else type_cast_2606_wire_constant;
    -- flow-through select operator MUX_2617_inst
    IMA14_2618 <= type_cast_2614_wire_constant when (BITSEL_u8_u1_2612_wire(0) /=  '0') else type_cast_2616_wire_constant;
    -- flow-through select operator MUX_2627_inst
    IMA15_2628 <= type_cast_2624_wire_constant when (BITSEL_u8_u1_2622_wire(0) /=  '0') else type_cast_2626_wire_constant;
    -- flow-through select operator MUX_2637_inst
    IMA16_2638 <= type_cast_2634_wire_constant when (BITSEL_u8_u1_2632_wire(0) /=  '0') else type_cast_2636_wire_constant;
    -- flow-through select operator MUX_2647_inst
    IMA17_2648 <= type_cast_2644_wire_constant when (BITSEL_u8_u1_2642_wire(0) /=  '0') else type_cast_2646_wire_constant;
    -- flow-through select operator MUX_2657_inst
    IMA18_2658 <= type_cast_2654_wire_constant when (BITSEL_u8_u1_2652_wire(0) /=  '0') else type_cast_2656_wire_constant;
    -- flow-through select operator MUX_2667_inst
    IMA19_2668 <= type_cast_2664_wire_constant when (BITSEL_u8_u1_2662_wire(0) /=  '0') else type_cast_2666_wire_constant;
    -- flow-through select operator MUX_2677_inst
    IMA20_2678 <= type_cast_2674_wire_constant when (BITSEL_u8_u1_2672_wire(0) /=  '0') else type_cast_2676_wire_constant;
    -- flow-through select operator MUX_2687_inst
    IMA21_2688 <= type_cast_2684_wire_constant when (BITSEL_u8_u1_2682_wire(0) /=  '0') else type_cast_2686_wire_constant;
    -- flow-through select operator MUX_2697_inst
    IMA22_2698 <= type_cast_2694_wire_constant when (BITSEL_u8_u1_2692_wire(0) /=  '0') else type_cast_2696_wire_constant;
    -- flow-through select operator MUX_2707_inst
    IMA23_2708 <= type_cast_2704_wire_constant when (BITSEL_u8_u1_2702_wire(0) /=  '0') else type_cast_2706_wire_constant;
    -- flow-through select operator MUX_2717_inst
    IMA24_2718 <= type_cast_2714_wire_constant when (BITSEL_u8_u1_2712_wire(0) /=  '0') else type_cast_2716_wire_constant;
    -- flow-through select operator MUX_2727_inst
    IMA25_2728 <= type_cast_2724_wire_constant when (BITSEL_u8_u1_2722_wire(0) /=  '0') else type_cast_2726_wire_constant;
    -- flow-through select operator MUX_2737_inst
    IMA26_2738 <= type_cast_2734_wire_constant when (BITSEL_u8_u1_2732_wire(0) /=  '0') else type_cast_2736_wire_constant;
    -- flow-through select operator MUX_2747_inst
    IMA27_2748 <= type_cast_2744_wire_constant when (BITSEL_u8_u1_2742_wire(0) /=  '0') else type_cast_2746_wire_constant;
    -- flow-through select operator MUX_2757_inst
    IMA28_2758 <= type_cast_2754_wire_constant when (BITSEL_u8_u1_2752_wire(0) /=  '0') else type_cast_2756_wire_constant;
    -- flow-through select operator MUX_2767_inst
    IMA29_2768 <= type_cast_2764_wire_constant when (BITSEL_u8_u1_2762_wire(0) /=  '0') else type_cast_2766_wire_constant;
    -- flow-through select operator MUX_2777_inst
    IMA30_2778 <= type_cast_2774_wire_constant when (BITSEL_u8_u1_2772_wire(0) /=  '0') else type_cast_2776_wire_constant;
    -- flow-through select operator MUX_2787_inst
    IMA31_2788 <= type_cast_2784_wire_constant when (BITSEL_u8_u1_2782_wire(0) /=  '0') else type_cast_2786_wire_constant;
    -- flow-through select operator MUX_2797_inst
    IMA32_2798 <= type_cast_2794_wire_constant when (BITSEL_u8_u1_2792_wire(0) /=  '0') else type_cast_2796_wire_constant;
    -- flow-through select operator MUX_2807_inst
    IMA33_2808 <= type_cast_2804_wire_constant when (BITSEL_u8_u1_2802_wire(0) /=  '0') else type_cast_2806_wire_constant;
    -- flow-through select operator MUX_2817_inst
    IMA34_2818 <= type_cast_2814_wire_constant when (BITSEL_u8_u1_2812_wire(0) /=  '0') else type_cast_2816_wire_constant;
    -- flow-through select operator MUX_2827_inst
    IMA35_2828 <= type_cast_2824_wire_constant when (BITSEL_u8_u1_2822_wire(0) /=  '0') else type_cast_2826_wire_constant;
    -- flow-through select operator MUX_2837_inst
    IMA36_2838 <= type_cast_2834_wire_constant when (BITSEL_u8_u1_2832_wire(0) /=  '0') else type_cast_2836_wire_constant;
    -- flow-through select operator MUX_2847_inst
    IMA37_2848 <= type_cast_2844_wire_constant when (BITSEL_u8_u1_2842_wire(0) /=  '0') else type_cast_2846_wire_constant;
    -- flow-through select operator MUX_2857_inst
    IMA38_2858 <= type_cast_2854_wire_constant when (BITSEL_u8_u1_2852_wire(0) /=  '0') else type_cast_2856_wire_constant;
    -- flow-through select operator MUX_2867_inst
    IMA39_2868 <= type_cast_2864_wire_constant when (BITSEL_u8_u1_2862_wire(0) /=  '0') else type_cast_2866_wire_constant;
    -- flow-through select operator MUX_2877_inst
    IMA40_2878 <= type_cast_2874_wire_constant when (BITSEL_u8_u1_2872_wire(0) /=  '0') else type_cast_2876_wire_constant;
    -- flow-through select operator MUX_2887_inst
    IMA41_2888 <= type_cast_2884_wire_constant when (BITSEL_u8_u1_2882_wire(0) /=  '0') else type_cast_2886_wire_constant;
    -- flow-through select operator MUX_2897_inst
    IMA42_2898 <= type_cast_2894_wire_constant when (BITSEL_u8_u1_2892_wire(0) /=  '0') else type_cast_2896_wire_constant;
    -- flow-through select operator MUX_2907_inst
    IMA43_2908 <= type_cast_2904_wire_constant when (BITSEL_u8_u1_2902_wire(0) /=  '0') else type_cast_2906_wire_constant;
    -- flow-through select operator MUX_2917_inst
    IMA44_2918 <= type_cast_2914_wire_constant when (BITSEL_u8_u1_2912_wire(0) /=  '0') else type_cast_2916_wire_constant;
    -- flow-through select operator MUX_2927_inst
    IMA45_2928 <= type_cast_2924_wire_constant when (BITSEL_u8_u1_2922_wire(0) /=  '0') else type_cast_2926_wire_constant;
    -- flow-through select operator MUX_2937_inst
    IMA46_2938 <= type_cast_2934_wire_constant when (BITSEL_u8_u1_2932_wire(0) /=  '0') else type_cast_2936_wire_constant;
    -- flow-through select operator MUX_2947_inst
    IMA47_2948 <= type_cast_2944_wire_constant when (BITSEL_u8_u1_2942_wire(0) /=  '0') else type_cast_2946_wire_constant;
    -- flow-through select operator MUX_2957_inst
    IMA48_2958 <= type_cast_2954_wire_constant when (BITSEL_u8_u1_2952_wire(0) /=  '0') else type_cast_2956_wire_constant;
    -- flow-through select operator MUX_2967_inst
    IMA49_2968 <= type_cast_2964_wire_constant when (BITSEL_u8_u1_2962_wire(0) /=  '0') else type_cast_2966_wire_constant;
    -- flow-through select operator MUX_2977_inst
    IMA50_2978 <= type_cast_2974_wire_constant when (BITSEL_u8_u1_2972_wire(0) /=  '0') else type_cast_2976_wire_constant;
    -- flow-through select operator MUX_2987_inst
    IMA51_2988 <= type_cast_2984_wire_constant when (BITSEL_u8_u1_2982_wire(0) /=  '0') else type_cast_2986_wire_constant;
    -- flow-through select operator MUX_2997_inst
    IMA52_2998 <= type_cast_2994_wire_constant when (BITSEL_u8_u1_2992_wire(0) /=  '0') else type_cast_2996_wire_constant;
    -- flow-through select operator MUX_3007_inst
    IMA53_3008 <= type_cast_3004_wire_constant when (BITSEL_u8_u1_3002_wire(0) /=  '0') else type_cast_3006_wire_constant;
    -- flow-through select operator MUX_3017_inst
    IMA54_3018 <= type_cast_3014_wire_constant when (BITSEL_u8_u1_3012_wire(0) /=  '0') else type_cast_3016_wire_constant;
    -- flow-through select operator MUX_3027_inst
    IMA55_3028 <= type_cast_3024_wire_constant when (BITSEL_u8_u1_3022_wire(0) /=  '0') else type_cast_3026_wire_constant;
    -- flow-through select operator MUX_3037_inst
    IMA56_3038 <= type_cast_3034_wire_constant when (BITSEL_u8_u1_3032_wire(0) /=  '0') else type_cast_3036_wire_constant;
    -- flow-through select operator MUX_3047_inst
    IMA57_3048 <= type_cast_3044_wire_constant when (BITSEL_u8_u1_3042_wire(0) /=  '0') else type_cast_3046_wire_constant;
    -- flow-through select operator MUX_3057_inst
    IMA58_3058 <= type_cast_3054_wire_constant when (BITSEL_u8_u1_3052_wire(0) /=  '0') else type_cast_3056_wire_constant;
    -- flow-through select operator MUX_3067_inst
    IMA59_3068 <= type_cast_3064_wire_constant when (BITSEL_u8_u1_3062_wire(0) /=  '0') else type_cast_3066_wire_constant;
    -- flow-through select operator MUX_3077_inst
    IMA60_3078 <= type_cast_3074_wire_constant when (BITSEL_u8_u1_3072_wire(0) /=  '0') else type_cast_3076_wire_constant;
    -- flow-through select operator MUX_3087_inst
    IMA61_3088 <= type_cast_3084_wire_constant when (BITSEL_u8_u1_3082_wire(0) /=  '0') else type_cast_3086_wire_constant;
    -- flow-through select operator MUX_3097_inst
    IMA62_3098 <= type_cast_3094_wire_constant when (BITSEL_u8_u1_3092_wire(0) /=  '0') else type_cast_3096_wire_constant;
    -- flow-through select operator MUX_3107_inst
    IMA63_3108 <= type_cast_3104_wire_constant when (BITSEL_u8_u1_3102_wire(0) /=  '0') else type_cast_3106_wire_constant;
    -- flow-through select operator MUX_3117_inst
    IMA64_3118 <= type_cast_3114_wire_constant when (BITSEL_u8_u1_3112_wire(0) /=  '0') else type_cast_3116_wire_constant;
    -- flow-through select operator MUX_3127_inst
    IMA65_3128 <= type_cast_3124_wire_constant when (BITSEL_u8_u1_3122_wire(0) /=  '0') else type_cast_3126_wire_constant;
    -- flow-through select operator MUX_3137_inst
    IMA66_3138 <= type_cast_3134_wire_constant when (BITSEL_u8_u1_3132_wire(0) /=  '0') else type_cast_3136_wire_constant;
    -- flow-through select operator MUX_3147_inst
    IMA67_3148 <= type_cast_3144_wire_constant when (BITSEL_u8_u1_3142_wire(0) /=  '0') else type_cast_3146_wire_constant;
    -- flow-through select operator MUX_3157_inst
    IMA68_3158 <= type_cast_3154_wire_constant when (BITSEL_u8_u1_3152_wire(0) /=  '0') else type_cast_3156_wire_constant;
    -- flow-through select operator MUX_3167_inst
    IMA69_3168 <= type_cast_3164_wire_constant when (BITSEL_u8_u1_3162_wire(0) /=  '0') else type_cast_3166_wire_constant;
    -- flow-through select operator MUX_3177_inst
    IMA70_3178 <= type_cast_3174_wire_constant when (BITSEL_u8_u1_3172_wire(0) /=  '0') else type_cast_3176_wire_constant;
    -- flow-through select operator MUX_3187_inst
    IMA71_3188 <= type_cast_3184_wire_constant when (BITSEL_u8_u1_3182_wire(0) /=  '0') else type_cast_3186_wire_constant;
    -- flow-through select operator MUX_3197_inst
    IMA72_3198 <= type_cast_3194_wire_constant when (BITSEL_u8_u1_3192_wire(0) /=  '0') else type_cast_3196_wire_constant;
    -- flow-through select operator MUX_3207_inst
    IMA73_3208 <= type_cast_3204_wire_constant when (BITSEL_u8_u1_3202_wire(0) /=  '0') else type_cast_3206_wire_constant;
    -- flow-through select operator MUX_3217_inst
    IMA74_3218 <= type_cast_3214_wire_constant when (BITSEL_u8_u1_3212_wire(0) /=  '0') else type_cast_3216_wire_constant;
    -- flow-through select operator MUX_3227_inst
    IMA75_3228 <= type_cast_3224_wire_constant when (BITSEL_u8_u1_3222_wire(0) /=  '0') else type_cast_3226_wire_constant;
    -- flow-through select operator MUX_3237_inst
    IMA76_3238 <= type_cast_3234_wire_constant when (BITSEL_u8_u1_3232_wire(0) /=  '0') else type_cast_3236_wire_constant;
    -- flow-through select operator MUX_3247_inst
    IMA77_3248 <= type_cast_3244_wire_constant when (BITSEL_u8_u1_3242_wire(0) /=  '0') else type_cast_3246_wire_constant;
    -- flow-through select operator MUX_3257_inst
    IMA78_3258 <= type_cast_3254_wire_constant when (BITSEL_u8_u1_3252_wire(0) /=  '0') else type_cast_3256_wire_constant;
    -- flow-through select operator MUX_3267_inst
    IMA79_3268 <= type_cast_3264_wire_constant when (BITSEL_u8_u1_3262_wire(0) /=  '0') else type_cast_3266_wire_constant;
    -- flow-through select operator MUX_3277_inst
    IMA80_3278 <= type_cast_3274_wire_constant when (BITSEL_u8_u1_3272_wire(0) /=  '0') else type_cast_3276_wire_constant;
    -- flow-through select operator MUX_3287_inst
    IMA81_3288 <= type_cast_3284_wire_constant when (BITSEL_u8_u1_3282_wire(0) /=  '0') else type_cast_3286_wire_constant;
    -- flow-through select operator MUX_3297_inst
    IMA82_3298 <= type_cast_3294_wire_constant when (BITSEL_u8_u1_3292_wire(0) /=  '0') else type_cast_3296_wire_constant;
    -- flow-through select operator MUX_3307_inst
    IMA83_3308 <= type_cast_3304_wire_constant when (BITSEL_u8_u1_3302_wire(0) /=  '0') else type_cast_3306_wire_constant;
    -- flow-through select operator MUX_3317_inst
    IMA84_3318 <= type_cast_3314_wire_constant when (BITSEL_u8_u1_3312_wire(0) /=  '0') else type_cast_3316_wire_constant;
    -- flow-through select operator MUX_3327_inst
    IMA85_3328 <= type_cast_3324_wire_constant when (BITSEL_u8_u1_3322_wire(0) /=  '0') else type_cast_3326_wire_constant;
    -- flow-through select operator MUX_3337_inst
    IMA86_3338 <= type_cast_3334_wire_constant when (BITSEL_u8_u1_3332_wire(0) /=  '0') else type_cast_3336_wire_constant;
    -- flow-through select operator MUX_3347_inst
    IMA87_3348 <= type_cast_3344_wire_constant when (BITSEL_u8_u1_3342_wire(0) /=  '0') else type_cast_3346_wire_constant;
    -- flow-through select operator MUX_3357_inst
    IMA88_3358 <= type_cast_3354_wire_constant when (BITSEL_u8_u1_3352_wire(0) /=  '0') else type_cast_3356_wire_constant;
    -- flow-through select operator MUX_3367_inst
    IMA89_3368 <= type_cast_3364_wire_constant when (BITSEL_u8_u1_3362_wire(0) /=  '0') else type_cast_3366_wire_constant;
    -- flow-through select operator MUX_3377_inst
    IMA90_3378 <= type_cast_3374_wire_constant when (BITSEL_u8_u1_3372_wire(0) /=  '0') else type_cast_3376_wire_constant;
    -- flow-through select operator MUX_3387_inst
    IMA91_3388 <= type_cast_3384_wire_constant when (BITSEL_u8_u1_3382_wire(0) /=  '0') else type_cast_3386_wire_constant;
    -- flow-through select operator MUX_3397_inst
    IMA92_3398 <= type_cast_3394_wire_constant when (BITSEL_u8_u1_3392_wire(0) /=  '0') else type_cast_3396_wire_constant;
    -- flow-through select operator MUX_3407_inst
    IMA93_3408 <= type_cast_3404_wire_constant when (BITSEL_u8_u1_3402_wire(0) /=  '0') else type_cast_3406_wire_constant;
    -- flow-through select operator MUX_3417_inst
    IMA94_3418 <= type_cast_3414_wire_constant when (BITSEL_u8_u1_3412_wire(0) /=  '0') else type_cast_3416_wire_constant;
    -- flow-through select operator MUX_3427_inst
    IMA95_3428 <= type_cast_3424_wire_constant when (BITSEL_u8_u1_3422_wire(0) /=  '0') else type_cast_3426_wire_constant;
    -- flow-through select operator MUX_3437_inst
    IMA96_3438 <= type_cast_3434_wire_constant when (BITSEL_u8_u1_3432_wire(0) /=  '0') else type_cast_3436_wire_constant;
    -- flow-through select operator MUX_3447_inst
    IMA97_3448 <= type_cast_3444_wire_constant when (BITSEL_u8_u1_3442_wire(0) /=  '0') else type_cast_3446_wire_constant;
    -- flow-through select operator MUX_3457_inst
    IMA98_3458 <= type_cast_3454_wire_constant when (BITSEL_u8_u1_3452_wire(0) /=  '0') else type_cast_3456_wire_constant;
    -- flow-through select operator MUX_3467_inst
    IMA99_3468 <= type_cast_3464_wire_constant when (BITSEL_u8_u1_3462_wire(0) /=  '0') else type_cast_3466_wire_constant;
    -- flow-through select operator MUX_3477_inst
    IMA100_3478 <= type_cast_3474_wire_constant when (BITSEL_u8_u1_3472_wire(0) /=  '0') else type_cast_3476_wire_constant;
    -- flow-through select operator MUX_3487_inst
    IMA101_3488 <= type_cast_3484_wire_constant when (BITSEL_u8_u1_3482_wire(0) /=  '0') else type_cast_3486_wire_constant;
    -- flow-through select operator MUX_3497_inst
    IMA102_3498 <= type_cast_3494_wire_constant when (BITSEL_u8_u1_3492_wire(0) /=  '0') else type_cast_3496_wire_constant;
    -- flow-through select operator MUX_3507_inst
    IMA103_3508 <= type_cast_3504_wire_constant when (BITSEL_u8_u1_3502_wire(0) /=  '0') else type_cast_3506_wire_constant;
    -- flow-through select operator MUX_3517_inst
    IMA104_3518 <= type_cast_3514_wire_constant when (BITSEL_u8_u1_3512_wire(0) /=  '0') else type_cast_3516_wire_constant;
    -- flow-through select operator MUX_3527_inst
    IMA105_3528 <= type_cast_3524_wire_constant when (BITSEL_u8_u1_3522_wire(0) /=  '0') else type_cast_3526_wire_constant;
    -- flow-through select operator MUX_3537_inst
    IMA106_3538 <= type_cast_3534_wire_constant when (BITSEL_u8_u1_3532_wire(0) /=  '0') else type_cast_3536_wire_constant;
    -- flow-through select operator MUX_3547_inst
    IMA107_3548 <= type_cast_3544_wire_constant when (BITSEL_u8_u1_3542_wire(0) /=  '0') else type_cast_3546_wire_constant;
    -- flow-through select operator MUX_3557_inst
    IMA108_3558 <= type_cast_3554_wire_constant when (BITSEL_u8_u1_3552_wire(0) /=  '0') else type_cast_3556_wire_constant;
    -- flow-through select operator MUX_3567_inst
    IMA109_3568 <= type_cast_3564_wire_constant when (BITSEL_u8_u1_3562_wire(0) /=  '0') else type_cast_3566_wire_constant;
    -- flow-through select operator MUX_3577_inst
    IMA110_3578 <= type_cast_3574_wire_constant when (BITSEL_u8_u1_3572_wire(0) /=  '0') else type_cast_3576_wire_constant;
    -- flow-through select operator MUX_3587_inst
    IMA111_3588 <= type_cast_3584_wire_constant when (BITSEL_u8_u1_3582_wire(0) /=  '0') else type_cast_3586_wire_constant;
    -- flow-through select operator MUX_3597_inst
    IMA112_3598 <= type_cast_3594_wire_constant when (BITSEL_u8_u1_3592_wire(0) /=  '0') else type_cast_3596_wire_constant;
    -- flow-through select operator MUX_3607_inst
    IMA113_3608 <= type_cast_3604_wire_constant when (BITSEL_u8_u1_3602_wire(0) /=  '0') else type_cast_3606_wire_constant;
    -- flow-through select operator MUX_3617_inst
    IMA114_3618 <= type_cast_3614_wire_constant when (BITSEL_u8_u1_3612_wire(0) /=  '0') else type_cast_3616_wire_constant;
    -- flow-through select operator MUX_3627_inst
    IMA115_3628 <= type_cast_3624_wire_constant when (BITSEL_u8_u1_3622_wire(0) /=  '0') else type_cast_3626_wire_constant;
    -- flow-through select operator MUX_3637_inst
    IMA116_3638 <= type_cast_3634_wire_constant when (BITSEL_u8_u1_3632_wire(0) /=  '0') else type_cast_3636_wire_constant;
    -- flow-through select operator MUX_3647_inst
    IMA117_3648 <= type_cast_3644_wire_constant when (BITSEL_u8_u1_3642_wire(0) /=  '0') else type_cast_3646_wire_constant;
    -- flow-through select operator MUX_3657_inst
    IMA118_3658 <= type_cast_3654_wire_constant when (BITSEL_u8_u1_3652_wire(0) /=  '0') else type_cast_3656_wire_constant;
    -- flow-through select operator MUX_3667_inst
    IMA119_3668 <= type_cast_3664_wire_constant when (BITSEL_u8_u1_3662_wire(0) /=  '0') else type_cast_3666_wire_constant;
    -- flow-through select operator MUX_3677_inst
    IMA120_3678 <= type_cast_3674_wire_constant when (BITSEL_u8_u1_3672_wire(0) /=  '0') else type_cast_3676_wire_constant;
    -- flow-through select operator MUX_3687_inst
    IMA121_3688 <= type_cast_3684_wire_constant when (BITSEL_u8_u1_3682_wire(0) /=  '0') else type_cast_3686_wire_constant;
    -- flow-through select operator MUX_3697_inst
    IMA122_3698 <= type_cast_3694_wire_constant when (BITSEL_u8_u1_3692_wire(0) /=  '0') else type_cast_3696_wire_constant;
    -- flow-through select operator MUX_3707_inst
    IMA123_3708 <= type_cast_3704_wire_constant when (BITSEL_u8_u1_3702_wire(0) /=  '0') else type_cast_3706_wire_constant;
    -- flow-through select operator MUX_3717_inst
    IMA124_3718 <= type_cast_3714_wire_constant when (BITSEL_u8_u1_3712_wire(0) /=  '0') else type_cast_3716_wire_constant;
    -- flow-through select operator MUX_3727_inst
    IMA125_3728 <= type_cast_3724_wire_constant when (BITSEL_u8_u1_3722_wire(0) /=  '0') else type_cast_3726_wire_constant;
    -- flow-through select operator MUX_3737_inst
    IMA126_3738 <= type_cast_3734_wire_constant when (BITSEL_u8_u1_3732_wire(0) /=  '0') else type_cast_3736_wire_constant;
    -- flow-through select operator MUX_3747_inst
    IMA127_3748 <= type_cast_3744_wire_constant when (BITSEL_u8_u1_3742_wire(0) /=  '0') else type_cast_3746_wire_constant;
    -- flow-through select operator MUX_3755_inst
    IMB0_3756 <= IMA1_2488 when (BITSEL_u8_u1_3752_wire(0) /=  '0') else IMA0_2478;
    -- flow-through select operator MUX_3763_inst
    IMB1_3764 <= IMA3_2508 when (BITSEL_u8_u1_3760_wire(0) /=  '0') else IMA2_2498;
    -- flow-through select operator MUX_3771_inst
    IMB2_3772 <= IMA5_2528 when (BITSEL_u8_u1_3768_wire(0) /=  '0') else IMA4_2518;
    -- flow-through select operator MUX_3779_inst
    IMB3_3780 <= IMA7_2548 when (BITSEL_u8_u1_3776_wire(0) /=  '0') else IMA6_2538;
    -- flow-through select operator MUX_3787_inst
    IMB4_3788 <= IMA9_2568 when (BITSEL_u8_u1_3784_wire(0) /=  '0') else IMA8_2558;
    -- flow-through select operator MUX_3795_inst
    IMB5_3796 <= IMA11_2588 when (BITSEL_u8_u1_3792_wire(0) /=  '0') else IMA10_2578;
    -- flow-through select operator MUX_3803_inst
    IMB6_3804 <= IMA13_2608 when (BITSEL_u8_u1_3800_wire(0) /=  '0') else IMA12_2598;
    -- flow-through select operator MUX_3811_inst
    IMB7_3812 <= IMA15_2628 when (BITSEL_u8_u1_3808_wire(0) /=  '0') else IMA14_2618;
    -- flow-through select operator MUX_3819_inst
    IMB8_3820 <= IMA17_2648 when (BITSEL_u8_u1_3816_wire(0) /=  '0') else IMA16_2638;
    -- flow-through select operator MUX_3827_inst
    IMB9_3828 <= IMA19_2668 when (BITSEL_u8_u1_3824_wire(0) /=  '0') else IMA18_2658;
    -- flow-through select operator MUX_3835_inst
    IMB10_3836 <= IMA21_2688 when (BITSEL_u8_u1_3832_wire(0) /=  '0') else IMA20_2678;
    -- flow-through select operator MUX_3843_inst
    IMB11_3844 <= IMA23_2708 when (BITSEL_u8_u1_3840_wire(0) /=  '0') else IMA22_2698;
    -- flow-through select operator MUX_3851_inst
    IMB12_3852 <= IMA25_2728 when (BITSEL_u8_u1_3848_wire(0) /=  '0') else IMA24_2718;
    -- flow-through select operator MUX_3859_inst
    IMB13_3860 <= IMA27_2748 when (BITSEL_u8_u1_3856_wire(0) /=  '0') else IMA26_2738;
    -- flow-through select operator MUX_3867_inst
    IMB14_3868 <= IMA29_2768 when (BITSEL_u8_u1_3864_wire(0) /=  '0') else IMA28_2758;
    -- flow-through select operator MUX_3875_inst
    IMB15_3876 <= IMA31_2788 when (BITSEL_u8_u1_3872_wire(0) /=  '0') else IMA30_2778;
    -- flow-through select operator MUX_3883_inst
    IMB16_3884 <= IMA33_2808 when (BITSEL_u8_u1_3880_wire(0) /=  '0') else IMA32_2798;
    -- flow-through select operator MUX_3891_inst
    IMB17_3892 <= IMA35_2828 when (BITSEL_u8_u1_3888_wire(0) /=  '0') else IMA34_2818;
    -- flow-through select operator MUX_3899_inst
    IMB18_3900 <= IMA37_2848 when (BITSEL_u8_u1_3896_wire(0) /=  '0') else IMA36_2838;
    -- flow-through select operator MUX_3907_inst
    IMB19_3908 <= IMA39_2868 when (BITSEL_u8_u1_3904_wire(0) /=  '0') else IMA38_2858;
    -- flow-through select operator MUX_3915_inst
    IMB20_3916 <= IMA41_2888 when (BITSEL_u8_u1_3912_wire(0) /=  '0') else IMA40_2878;
    -- flow-through select operator MUX_3923_inst
    IMB21_3924 <= IMA43_2908 when (BITSEL_u8_u1_3920_wire(0) /=  '0') else IMA42_2898;
    -- flow-through select operator MUX_3931_inst
    IMB22_3932 <= IMA45_2928 when (BITSEL_u8_u1_3928_wire(0) /=  '0') else IMA44_2918;
    -- flow-through select operator MUX_3939_inst
    IMB23_3940 <= IMA47_2948 when (BITSEL_u8_u1_3936_wire(0) /=  '0') else IMA46_2938;
    -- flow-through select operator MUX_3947_inst
    IMB24_3948 <= IMA49_2968 when (BITSEL_u8_u1_3944_wire(0) /=  '0') else IMA48_2958;
    -- flow-through select operator MUX_3955_inst
    IMB25_3956 <= IMA51_2988 when (BITSEL_u8_u1_3952_wire(0) /=  '0') else IMA50_2978;
    -- flow-through select operator MUX_3963_inst
    IMB26_3964 <= IMA53_3008 when (BITSEL_u8_u1_3960_wire(0) /=  '0') else IMA52_2998;
    -- flow-through select operator MUX_3971_inst
    IMB27_3972 <= IMA55_3028 when (BITSEL_u8_u1_3968_wire(0) /=  '0') else IMA54_3018;
    -- flow-through select operator MUX_3979_inst
    IMB28_3980 <= IMA57_3048 when (BITSEL_u8_u1_3976_wire(0) /=  '0') else IMA56_3038;
    -- flow-through select operator MUX_3987_inst
    IMB29_3988 <= IMA59_3068 when (BITSEL_u8_u1_3984_wire(0) /=  '0') else IMA58_3058;
    -- flow-through select operator MUX_3995_inst
    IMB30_3996 <= IMA61_3088 when (BITSEL_u8_u1_3992_wire(0) /=  '0') else IMA60_3078;
    -- flow-through select operator MUX_4003_inst
    IMB31_4004 <= IMA63_3108 when (BITSEL_u8_u1_4000_wire(0) /=  '0') else IMA62_3098;
    -- flow-through select operator MUX_4011_inst
    IMB32_4012 <= IMA65_3128 when (BITSEL_u8_u1_4008_wire(0) /=  '0') else IMA64_3118;
    -- flow-through select operator MUX_4019_inst
    IMB33_4020 <= IMA67_3148 when (BITSEL_u8_u1_4016_wire(0) /=  '0') else IMA66_3138;
    -- flow-through select operator MUX_4027_inst
    IMB34_4028 <= IMA69_3168 when (BITSEL_u8_u1_4024_wire(0) /=  '0') else IMA68_3158;
    -- flow-through select operator MUX_4035_inst
    IMB35_4036 <= IMA71_3188 when (BITSEL_u8_u1_4032_wire(0) /=  '0') else IMA70_3178;
    -- flow-through select operator MUX_4043_inst
    IMB36_4044 <= IMA73_3208 when (BITSEL_u8_u1_4040_wire(0) /=  '0') else IMA72_3198;
    -- flow-through select operator MUX_4051_inst
    IMB37_4052 <= IMA75_3228 when (BITSEL_u8_u1_4048_wire(0) /=  '0') else IMA74_3218;
    -- flow-through select operator MUX_4059_inst
    IMB38_4060 <= IMA77_3248 when (BITSEL_u8_u1_4056_wire(0) /=  '0') else IMA76_3238;
    -- flow-through select operator MUX_4067_inst
    IMB39_4068 <= IMA79_3268 when (BITSEL_u8_u1_4064_wire(0) /=  '0') else IMA78_3258;
    -- flow-through select operator MUX_4075_inst
    IMB40_4076 <= IMA81_3288 when (BITSEL_u8_u1_4072_wire(0) /=  '0') else IMA80_3278;
    -- flow-through select operator MUX_4083_inst
    IMB41_4084 <= IMA83_3308 when (BITSEL_u8_u1_4080_wire(0) /=  '0') else IMA82_3298;
    -- flow-through select operator MUX_4091_inst
    IMB42_4092 <= IMA85_3328 when (BITSEL_u8_u1_4088_wire(0) /=  '0') else IMA84_3318;
    -- flow-through select operator MUX_4099_inst
    IMB43_4100 <= IMA87_3348 when (BITSEL_u8_u1_4096_wire(0) /=  '0') else IMA86_3338;
    -- flow-through select operator MUX_4107_inst
    IMB44_4108 <= IMA89_3368 when (BITSEL_u8_u1_4104_wire(0) /=  '0') else IMA88_3358;
    -- flow-through select operator MUX_4115_inst
    IMB45_4116 <= IMA91_3388 when (BITSEL_u8_u1_4112_wire(0) /=  '0') else IMA90_3378;
    -- flow-through select operator MUX_4123_inst
    IMB46_4124 <= IMA93_3408 when (BITSEL_u8_u1_4120_wire(0) /=  '0') else IMA92_3398;
    -- flow-through select operator MUX_4131_inst
    IMB47_4132 <= IMA95_3428 when (BITSEL_u8_u1_4128_wire(0) /=  '0') else IMA94_3418;
    -- flow-through select operator MUX_4139_inst
    IMB48_4140 <= IMA97_3448 when (BITSEL_u8_u1_4136_wire(0) /=  '0') else IMA96_3438;
    -- flow-through select operator MUX_4147_inst
    IMB49_4148 <= IMA99_3468 when (BITSEL_u8_u1_4144_wire(0) /=  '0') else IMA98_3458;
    -- flow-through select operator MUX_4155_inst
    IMB50_4156 <= IMA101_3488 when (BITSEL_u8_u1_4152_wire(0) /=  '0') else IMA100_3478;
    -- flow-through select operator MUX_4163_inst
    IMB51_4164 <= IMA103_3508 when (BITSEL_u8_u1_4160_wire(0) /=  '0') else IMA102_3498;
    -- flow-through select operator MUX_4171_inst
    IMB52_4172 <= IMA105_3528 when (BITSEL_u8_u1_4168_wire(0) /=  '0') else IMA104_3518;
    -- flow-through select operator MUX_4179_inst
    IMB53_4180 <= IMA107_3548 when (BITSEL_u8_u1_4176_wire(0) /=  '0') else IMA106_3538;
    -- flow-through select operator MUX_4187_inst
    IMB54_4188 <= IMA109_3568 when (BITSEL_u8_u1_4184_wire(0) /=  '0') else IMA108_3558;
    -- flow-through select operator MUX_4195_inst
    IMB55_4196 <= IMA111_3588 when (BITSEL_u8_u1_4192_wire(0) /=  '0') else IMA110_3578;
    -- flow-through select operator MUX_4203_inst
    IMB56_4204 <= IMA113_3608 when (BITSEL_u8_u1_4200_wire(0) /=  '0') else IMA112_3598;
    -- flow-through select operator MUX_4211_inst
    IMB57_4212 <= IMA115_3628 when (BITSEL_u8_u1_4208_wire(0) /=  '0') else IMA114_3618;
    -- flow-through select operator MUX_4219_inst
    IMB58_4220 <= IMA117_3648 when (BITSEL_u8_u1_4216_wire(0) /=  '0') else IMA116_3638;
    -- flow-through select operator MUX_4227_inst
    IMB59_4228 <= IMA119_3668 when (BITSEL_u8_u1_4224_wire(0) /=  '0') else IMA118_3658;
    -- flow-through select operator MUX_4235_inst
    IMB60_4236 <= IMA121_3688 when (BITSEL_u8_u1_4232_wire(0) /=  '0') else IMA120_3678;
    -- flow-through select operator MUX_4243_inst
    IMB61_4244 <= IMA123_3708 when (BITSEL_u8_u1_4240_wire(0) /=  '0') else IMA122_3698;
    -- flow-through select operator MUX_4251_inst
    IMB62_4252 <= IMA125_3728 when (BITSEL_u8_u1_4248_wire(0) /=  '0') else IMA124_3718;
    -- flow-through select operator MUX_4259_inst
    IMB63_4260 <= IMA127_3748 when (BITSEL_u8_u1_4256_wire(0) /=  '0') else IMA126_3738;
    -- flow-through select operator MUX_4267_inst
    IMC0_4268 <= IMB1_3764 when (BITSEL_u8_u1_4264_wire(0) /=  '0') else IMB0_3756;
    -- flow-through select operator MUX_4275_inst
    IMC1_4276 <= IMB3_3780 when (BITSEL_u8_u1_4272_wire(0) /=  '0') else IMB2_3772;
    -- flow-through select operator MUX_4283_inst
    IMC2_4284 <= IMB5_3796 when (BITSEL_u8_u1_4280_wire(0) /=  '0') else IMB4_3788;
    -- flow-through select operator MUX_4291_inst
    IMC3_4292 <= IMB7_3812 when (BITSEL_u8_u1_4288_wire(0) /=  '0') else IMB6_3804;
    -- flow-through select operator MUX_4299_inst
    IMC4_4300 <= IMB9_3828 when (BITSEL_u8_u1_4296_wire(0) /=  '0') else IMB8_3820;
    -- flow-through select operator MUX_4307_inst
    IMC5_4308 <= IMB11_3844 when (BITSEL_u8_u1_4304_wire(0) /=  '0') else IMB10_3836;
    -- flow-through select operator MUX_4315_inst
    IMC6_4316 <= IMB13_3860 when (BITSEL_u8_u1_4312_wire(0) /=  '0') else IMB12_3852;
    -- flow-through select operator MUX_4323_inst
    IMC7_4324 <= IMB15_3876 when (BITSEL_u8_u1_4320_wire(0) /=  '0') else IMB14_3868;
    -- flow-through select operator MUX_4331_inst
    IMC8_4332 <= IMB17_3892 when (BITSEL_u8_u1_4328_wire(0) /=  '0') else IMB16_3884;
    -- flow-through select operator MUX_4339_inst
    IMC9_4340 <= IMB19_3908 when (BITSEL_u8_u1_4336_wire(0) /=  '0') else IMB18_3900;
    -- flow-through select operator MUX_4347_inst
    IMC10_4348 <= IMB21_3924 when (BITSEL_u8_u1_4344_wire(0) /=  '0') else IMB20_3916;
    -- flow-through select operator MUX_4355_inst
    IMC11_4356 <= IMB23_3940 when (BITSEL_u8_u1_4352_wire(0) /=  '0') else IMB22_3932;
    -- flow-through select operator MUX_4363_inst
    IMC12_4364 <= IMB25_3956 when (BITSEL_u8_u1_4360_wire(0) /=  '0') else IMB24_3948;
    -- flow-through select operator MUX_4371_inst
    IMC13_4372 <= IMB27_3972 when (BITSEL_u8_u1_4368_wire(0) /=  '0') else IMB26_3964;
    -- flow-through select operator MUX_4379_inst
    IMC14_4380 <= IMB29_3988 when (BITSEL_u8_u1_4376_wire(0) /=  '0') else IMB28_3980;
    -- flow-through select operator MUX_4387_inst
    IMC15_4388 <= IMB31_4004 when (BITSEL_u8_u1_4384_wire(0) /=  '0') else IMB30_3996;
    -- flow-through select operator MUX_4395_inst
    IMC16_4396 <= IMB33_4020 when (BITSEL_u8_u1_4392_wire(0) /=  '0') else IMB32_4012;
    -- flow-through select operator MUX_4403_inst
    IMC17_4404 <= IMB35_4036 when (BITSEL_u8_u1_4400_wire(0) /=  '0') else IMB34_4028;
    -- flow-through select operator MUX_4411_inst
    IMC18_4412 <= IMB37_4052 when (BITSEL_u8_u1_4408_wire(0) /=  '0') else IMB36_4044;
    -- flow-through select operator MUX_4419_inst
    IMC19_4420 <= IMB39_4068 when (BITSEL_u8_u1_4416_wire(0) /=  '0') else IMB38_4060;
    -- flow-through select operator MUX_4427_inst
    IMC20_4428 <= IMB41_4084 when (BITSEL_u8_u1_4424_wire(0) /=  '0') else IMB40_4076;
    -- flow-through select operator MUX_4435_inst
    IMC21_4436 <= IMB43_4100 when (BITSEL_u8_u1_4432_wire(0) /=  '0') else IMB42_4092;
    -- flow-through select operator MUX_4443_inst
    IMC22_4444 <= IMB45_4116 when (BITSEL_u8_u1_4440_wire(0) /=  '0') else IMB44_4108;
    -- flow-through select operator MUX_4451_inst
    IMC23_4452 <= IMB47_4132 when (BITSEL_u8_u1_4448_wire(0) /=  '0') else IMB46_4124;
    -- flow-through select operator MUX_4459_inst
    IMC24_4460 <= IMB49_4148 when (BITSEL_u8_u1_4456_wire(0) /=  '0') else IMB48_4140;
    -- flow-through select operator MUX_4467_inst
    IMC25_4468 <= IMB51_4164 when (BITSEL_u8_u1_4464_wire(0) /=  '0') else IMB50_4156;
    -- flow-through select operator MUX_4475_inst
    IMC26_4476 <= IMB53_4180 when (BITSEL_u8_u1_4472_wire(0) /=  '0') else IMB52_4172;
    -- flow-through select operator MUX_4483_inst
    IMC27_4484 <= IMB55_4196 when (BITSEL_u8_u1_4480_wire(0) /=  '0') else IMB54_4188;
    -- flow-through select operator MUX_4491_inst
    IMC28_4492 <= IMB57_4212 when (BITSEL_u8_u1_4488_wire(0) /=  '0') else IMB56_4204;
    -- flow-through select operator MUX_4499_inst
    IMC29_4500 <= IMB59_4228 when (BITSEL_u8_u1_4496_wire(0) /=  '0') else IMB58_4220;
    -- flow-through select operator MUX_4507_inst
    IMC30_4508 <= IMB61_4244 when (BITSEL_u8_u1_4504_wire(0) /=  '0') else IMB60_4236;
    -- flow-through select operator MUX_4515_inst
    IMC31_4516 <= IMB63_4260 when (BITSEL_u8_u1_4512_wire(0) /=  '0') else IMB62_4252;
    -- flow-through select operator MUX_4523_inst
    IMD0_4524 <= IMC1_4276 when (BITSEL_u8_u1_4520_wire(0) /=  '0') else IMC0_4268;
    -- flow-through select operator MUX_4531_inst
    IMD1_4532 <= IMC3_4292 when (BITSEL_u8_u1_4528_wire(0) /=  '0') else IMC2_4284;
    -- flow-through select operator MUX_4539_inst
    IMD2_4540 <= IMC5_4308 when (BITSEL_u8_u1_4536_wire(0) /=  '0') else IMC4_4300;
    -- flow-through select operator MUX_4547_inst
    IMD3_4548 <= IMC7_4324 when (BITSEL_u8_u1_4544_wire(0) /=  '0') else IMC6_4316;
    -- flow-through select operator MUX_4555_inst
    IMD4_4556 <= IMC9_4340 when (BITSEL_u8_u1_4552_wire(0) /=  '0') else IMC8_4332;
    -- flow-through select operator MUX_4563_inst
    IMD5_4564 <= IMC11_4356 when (BITSEL_u8_u1_4560_wire(0) /=  '0') else IMC10_4348;
    -- flow-through select operator MUX_4571_inst
    IMD6_4572 <= IMC13_4372 when (BITSEL_u8_u1_4568_wire(0) /=  '0') else IMC12_4364;
    -- flow-through select operator MUX_4579_inst
    IMD7_4580 <= IMC15_4388 when (BITSEL_u8_u1_4576_wire(0) /=  '0') else IMC14_4380;
    -- flow-through select operator MUX_4587_inst
    IMD8_4588 <= IMC17_4404 when (BITSEL_u8_u1_4584_wire(0) /=  '0') else IMC16_4396;
    -- flow-through select operator MUX_4595_inst
    IMD9_4596 <= IMC19_4420 when (BITSEL_u8_u1_4592_wire(0) /=  '0') else IMC18_4412;
    -- flow-through select operator MUX_4603_inst
    IMD10_4604 <= IMC21_4436 when (BITSEL_u8_u1_4600_wire(0) /=  '0') else IMC20_4428;
    -- flow-through select operator MUX_4611_inst
    IMD11_4612 <= IMC23_4452 when (BITSEL_u8_u1_4608_wire(0) /=  '0') else IMC22_4444;
    -- flow-through select operator MUX_4619_inst
    IMD12_4620 <= IMC25_4468 when (BITSEL_u8_u1_4616_wire(0) /=  '0') else IMC24_4460;
    -- flow-through select operator MUX_4627_inst
    IMD13_4628 <= IMC27_4484 when (BITSEL_u8_u1_4624_wire(0) /=  '0') else IMC26_4476;
    -- flow-through select operator MUX_4635_inst
    IMD14_4636 <= IMC29_4500 when (BITSEL_u8_u1_4632_wire(0) /=  '0') else IMC28_4492;
    -- flow-through select operator MUX_4643_inst
    IMD15_4644 <= IMC31_4516 when (BITSEL_u8_u1_4640_wire(0) /=  '0') else IMC30_4508;
    -- flow-through select operator MUX_4651_inst
    IME0_4652 <= IMD1_4532 when (BITSEL_u8_u1_4648_wire(0) /=  '0') else IMD0_4524;
    -- flow-through select operator MUX_4659_inst
    IME1_4660 <= IMD3_4548 when (BITSEL_u8_u1_4656_wire(0) /=  '0') else IMD2_4540;
    -- flow-through select operator MUX_4667_inst
    IME2_4668 <= IMD5_4564 when (BITSEL_u8_u1_4664_wire(0) /=  '0') else IMD4_4556;
    -- flow-through select operator MUX_4675_inst
    IME3_4676 <= IMD7_4580 when (BITSEL_u8_u1_4672_wire(0) /=  '0') else IMD6_4572;
    -- flow-through select operator MUX_4683_inst
    IME4_4684 <= IMD9_4596 when (BITSEL_u8_u1_4680_wire(0) /=  '0') else IMD8_4588;
    -- flow-through select operator MUX_4691_inst
    IME5_4692 <= IMD11_4612 when (BITSEL_u8_u1_4688_wire(0) /=  '0') else IMD10_4604;
    -- flow-through select operator MUX_4699_inst
    IME6_4700 <= IMD13_4628 when (BITSEL_u8_u1_4696_wire(0) /=  '0') else IMD12_4620;
    -- flow-through select operator MUX_4707_inst
    IME7_4708 <= IMD15_4644 when (BITSEL_u8_u1_4704_wire(0) /=  '0') else IMD14_4636;
    -- flow-through select operator MUX_4715_inst
    IMF0_4716 <= IME1_4660 when (BITSEL_u8_u1_4712_wire(0) /=  '0') else IME0_4652;
    -- flow-through select operator MUX_4723_inst
    IMF1_4724 <= IME3_4676 when (BITSEL_u8_u1_4720_wire(0) /=  '0') else IME2_4668;
    -- flow-through select operator MUX_4731_inst
    IMF2_4732 <= IME5_4692 when (BITSEL_u8_u1_4728_wire(0) /=  '0') else IME4_4684;
    -- flow-through select operator MUX_4739_inst
    IMF3_4740 <= IME7_4708 when (BITSEL_u8_u1_4736_wire(0) /=  '0') else IME6_4700;
    -- flow-through select operator MUX_4747_inst
    IMG0_4748 <= IMF1_4724 when (BITSEL_u8_u1_4744_wire(0) /=  '0') else IMF0_4716;
    -- flow-through select operator MUX_4755_inst
    IMG1_4756 <= IMF3_4740 when (BITSEL_u8_u1_4752_wire(0) /=  '0') else IMF2_4732;
    -- flow-through select operator MUX_4763_inst
    s_out_buffer <= IMG1_4756 when (BITSEL_u8_u1_4760_wire(0) /=  '0') else IMG0_4748;
    -- binary operator BITSEL_u8_u1_2472_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2471_wire_constant, tmp_var);
      BITSEL_u8_u1_2472_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2482_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2481_wire_constant, tmp_var);
      BITSEL_u8_u1_2482_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2492_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2491_wire_constant, tmp_var);
      BITSEL_u8_u1_2492_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2502_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2501_wire_constant, tmp_var);
      BITSEL_u8_u1_2502_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2512_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2511_wire_constant, tmp_var);
      BITSEL_u8_u1_2512_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2522_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2521_wire_constant, tmp_var);
      BITSEL_u8_u1_2522_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2532_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2531_wire_constant, tmp_var);
      BITSEL_u8_u1_2532_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2542_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2541_wire_constant, tmp_var);
      BITSEL_u8_u1_2542_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2552_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2551_wire_constant, tmp_var);
      BITSEL_u8_u1_2552_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2562_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2561_wire_constant, tmp_var);
      BITSEL_u8_u1_2562_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2572_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2571_wire_constant, tmp_var);
      BITSEL_u8_u1_2572_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2582_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2581_wire_constant, tmp_var);
      BITSEL_u8_u1_2582_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2592_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2591_wire_constant, tmp_var);
      BITSEL_u8_u1_2592_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2602_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2601_wire_constant, tmp_var);
      BITSEL_u8_u1_2602_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2612_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2611_wire_constant, tmp_var);
      BITSEL_u8_u1_2612_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2622_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2621_wire_constant, tmp_var);
      BITSEL_u8_u1_2622_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2632_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2631_wire_constant, tmp_var);
      BITSEL_u8_u1_2632_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2642_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2641_wire_constant, tmp_var);
      BITSEL_u8_u1_2642_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2652_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2651_wire_constant, tmp_var);
      BITSEL_u8_u1_2652_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2662_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2661_wire_constant, tmp_var);
      BITSEL_u8_u1_2662_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2672_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2671_wire_constant, tmp_var);
      BITSEL_u8_u1_2672_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2682_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2681_wire_constant, tmp_var);
      BITSEL_u8_u1_2682_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2692_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2691_wire_constant, tmp_var);
      BITSEL_u8_u1_2692_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2702_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2701_wire_constant, tmp_var);
      BITSEL_u8_u1_2702_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2712_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2711_wire_constant, tmp_var);
      BITSEL_u8_u1_2712_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2722_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2721_wire_constant, tmp_var);
      BITSEL_u8_u1_2722_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2732_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2731_wire_constant, tmp_var);
      BITSEL_u8_u1_2732_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2742_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2741_wire_constant, tmp_var);
      BITSEL_u8_u1_2742_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2752_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2751_wire_constant, tmp_var);
      BITSEL_u8_u1_2752_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2762_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2761_wire_constant, tmp_var);
      BITSEL_u8_u1_2762_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2772_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2771_wire_constant, tmp_var);
      BITSEL_u8_u1_2772_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2782_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2781_wire_constant, tmp_var);
      BITSEL_u8_u1_2782_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2792_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2791_wire_constant, tmp_var);
      BITSEL_u8_u1_2792_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2802_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2801_wire_constant, tmp_var);
      BITSEL_u8_u1_2802_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2812_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2811_wire_constant, tmp_var);
      BITSEL_u8_u1_2812_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2822_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2821_wire_constant, tmp_var);
      BITSEL_u8_u1_2822_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2832_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2831_wire_constant, tmp_var);
      BITSEL_u8_u1_2832_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2842_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2841_wire_constant, tmp_var);
      BITSEL_u8_u1_2842_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2852_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2851_wire_constant, tmp_var);
      BITSEL_u8_u1_2852_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2862_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2861_wire_constant, tmp_var);
      BITSEL_u8_u1_2862_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2872_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2871_wire_constant, tmp_var);
      BITSEL_u8_u1_2872_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2882_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2881_wire_constant, tmp_var);
      BITSEL_u8_u1_2882_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2892_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2891_wire_constant, tmp_var);
      BITSEL_u8_u1_2892_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2902_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2901_wire_constant, tmp_var);
      BITSEL_u8_u1_2902_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2912_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2911_wire_constant, tmp_var);
      BITSEL_u8_u1_2912_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2922_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2921_wire_constant, tmp_var);
      BITSEL_u8_u1_2922_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2932_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2931_wire_constant, tmp_var);
      BITSEL_u8_u1_2932_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2942_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2941_wire_constant, tmp_var);
      BITSEL_u8_u1_2942_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2952_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2951_wire_constant, tmp_var);
      BITSEL_u8_u1_2952_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2962_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2961_wire_constant, tmp_var);
      BITSEL_u8_u1_2962_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2972_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2971_wire_constant, tmp_var);
      BITSEL_u8_u1_2972_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2982_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2981_wire_constant, tmp_var);
      BITSEL_u8_u1_2982_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_2992_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_2991_wire_constant, tmp_var);
      BITSEL_u8_u1_2992_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_3002_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3001_wire_constant, tmp_var);
      BITSEL_u8_u1_3002_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_3012_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3011_wire_constant, tmp_var);
      BITSEL_u8_u1_3012_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_3022_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3021_wire_constant, tmp_var);
      BITSEL_u8_u1_3022_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_3032_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3031_wire_constant, tmp_var);
      BITSEL_u8_u1_3032_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_3042_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3041_wire_constant, tmp_var);
      BITSEL_u8_u1_3042_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_3052_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3051_wire_constant, tmp_var);
      BITSEL_u8_u1_3052_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_3062_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3061_wire_constant, tmp_var);
      BITSEL_u8_u1_3062_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_3072_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3071_wire_constant, tmp_var);
      BITSEL_u8_u1_3072_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_3082_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3081_wire_constant, tmp_var);
      BITSEL_u8_u1_3082_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_3092_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3091_wire_constant, tmp_var);
      BITSEL_u8_u1_3092_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_3102_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3101_wire_constant, tmp_var);
      BITSEL_u8_u1_3102_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_3112_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3111_wire_constant, tmp_var);
      BITSEL_u8_u1_3112_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_3122_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3121_wire_constant, tmp_var);
      BITSEL_u8_u1_3122_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_3132_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3131_wire_constant, tmp_var);
      BITSEL_u8_u1_3132_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_3142_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3141_wire_constant, tmp_var);
      BITSEL_u8_u1_3142_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_3152_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3151_wire_constant, tmp_var);
      BITSEL_u8_u1_3152_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_3162_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3161_wire_constant, tmp_var);
      BITSEL_u8_u1_3162_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_3172_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3171_wire_constant, tmp_var);
      BITSEL_u8_u1_3172_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_3182_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3181_wire_constant, tmp_var);
      BITSEL_u8_u1_3182_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_3192_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3191_wire_constant, tmp_var);
      BITSEL_u8_u1_3192_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_3202_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3201_wire_constant, tmp_var);
      BITSEL_u8_u1_3202_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_3212_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3211_wire_constant, tmp_var);
      BITSEL_u8_u1_3212_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_3222_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3221_wire_constant, tmp_var);
      BITSEL_u8_u1_3222_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_3232_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3231_wire_constant, tmp_var);
      BITSEL_u8_u1_3232_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_3242_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3241_wire_constant, tmp_var);
      BITSEL_u8_u1_3242_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_3252_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3251_wire_constant, tmp_var);
      BITSEL_u8_u1_3252_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_3262_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3261_wire_constant, tmp_var);
      BITSEL_u8_u1_3262_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_3272_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3271_wire_constant, tmp_var);
      BITSEL_u8_u1_3272_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_3282_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3281_wire_constant, tmp_var);
      BITSEL_u8_u1_3282_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_3292_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3291_wire_constant, tmp_var);
      BITSEL_u8_u1_3292_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_3302_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3301_wire_constant, tmp_var);
      BITSEL_u8_u1_3302_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_3312_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3311_wire_constant, tmp_var);
      BITSEL_u8_u1_3312_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_3322_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3321_wire_constant, tmp_var);
      BITSEL_u8_u1_3322_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_3332_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3331_wire_constant, tmp_var);
      BITSEL_u8_u1_3332_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_3342_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3341_wire_constant, tmp_var);
      BITSEL_u8_u1_3342_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_3352_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3351_wire_constant, tmp_var);
      BITSEL_u8_u1_3352_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_3362_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3361_wire_constant, tmp_var);
      BITSEL_u8_u1_3362_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_3372_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3371_wire_constant, tmp_var);
      BITSEL_u8_u1_3372_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_3382_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3381_wire_constant, tmp_var);
      BITSEL_u8_u1_3382_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_3392_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3391_wire_constant, tmp_var);
      BITSEL_u8_u1_3392_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_3402_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3401_wire_constant, tmp_var);
      BITSEL_u8_u1_3402_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_3412_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3411_wire_constant, tmp_var);
      BITSEL_u8_u1_3412_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_3422_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3421_wire_constant, tmp_var);
      BITSEL_u8_u1_3422_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_3432_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3431_wire_constant, tmp_var);
      BITSEL_u8_u1_3432_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_3442_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3441_wire_constant, tmp_var);
      BITSEL_u8_u1_3442_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_3452_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3451_wire_constant, tmp_var);
      BITSEL_u8_u1_3452_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_3462_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3461_wire_constant, tmp_var);
      BITSEL_u8_u1_3462_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_3472_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3471_wire_constant, tmp_var);
      BITSEL_u8_u1_3472_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_3482_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3481_wire_constant, tmp_var);
      BITSEL_u8_u1_3482_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_3492_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3491_wire_constant, tmp_var);
      BITSEL_u8_u1_3492_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_3502_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3501_wire_constant, tmp_var);
      BITSEL_u8_u1_3502_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_3512_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3511_wire_constant, tmp_var);
      BITSEL_u8_u1_3512_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_3522_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3521_wire_constant, tmp_var);
      BITSEL_u8_u1_3522_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_3532_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3531_wire_constant, tmp_var);
      BITSEL_u8_u1_3532_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_3542_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3541_wire_constant, tmp_var);
      BITSEL_u8_u1_3542_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_3552_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3551_wire_constant, tmp_var);
      BITSEL_u8_u1_3552_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_3562_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3561_wire_constant, tmp_var);
      BITSEL_u8_u1_3562_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_3572_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3571_wire_constant, tmp_var);
      BITSEL_u8_u1_3572_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_3582_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3581_wire_constant, tmp_var);
      BITSEL_u8_u1_3582_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_3592_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3591_wire_constant, tmp_var);
      BITSEL_u8_u1_3592_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_3602_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3601_wire_constant, tmp_var);
      BITSEL_u8_u1_3602_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_3612_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3611_wire_constant, tmp_var);
      BITSEL_u8_u1_3612_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_3622_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3621_wire_constant, tmp_var);
      BITSEL_u8_u1_3622_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_3632_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3631_wire_constant, tmp_var);
      BITSEL_u8_u1_3632_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_3642_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3641_wire_constant, tmp_var);
      BITSEL_u8_u1_3642_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_3652_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3651_wire_constant, tmp_var);
      BITSEL_u8_u1_3652_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_3662_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3661_wire_constant, tmp_var);
      BITSEL_u8_u1_3662_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_3672_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3671_wire_constant, tmp_var);
      BITSEL_u8_u1_3672_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_3682_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3681_wire_constant, tmp_var);
      BITSEL_u8_u1_3682_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_3692_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3691_wire_constant, tmp_var);
      BITSEL_u8_u1_3692_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_3702_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3701_wire_constant, tmp_var);
      BITSEL_u8_u1_3702_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_3712_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3711_wire_constant, tmp_var);
      BITSEL_u8_u1_3712_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_3722_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3721_wire_constant, tmp_var);
      BITSEL_u8_u1_3722_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_3732_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3731_wire_constant, tmp_var);
      BITSEL_u8_u1_3732_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_3742_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3741_wire_constant, tmp_var);
      BITSEL_u8_u1_3742_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_3752_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3751_wire_constant, tmp_var);
      BITSEL_u8_u1_3752_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_3760_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3759_wire_constant, tmp_var);
      BITSEL_u8_u1_3760_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_3768_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3767_wire_constant, tmp_var);
      BITSEL_u8_u1_3768_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_3776_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3775_wire_constant, tmp_var);
      BITSEL_u8_u1_3776_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_3784_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3783_wire_constant, tmp_var);
      BITSEL_u8_u1_3784_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_3792_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3791_wire_constant, tmp_var);
      BITSEL_u8_u1_3792_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_3800_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3799_wire_constant, tmp_var);
      BITSEL_u8_u1_3800_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_3808_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3807_wire_constant, tmp_var);
      BITSEL_u8_u1_3808_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_3816_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3815_wire_constant, tmp_var);
      BITSEL_u8_u1_3816_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_3824_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3823_wire_constant, tmp_var);
      BITSEL_u8_u1_3824_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_3832_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3831_wire_constant, tmp_var);
      BITSEL_u8_u1_3832_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_3840_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3839_wire_constant, tmp_var);
      BITSEL_u8_u1_3840_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_3848_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3847_wire_constant, tmp_var);
      BITSEL_u8_u1_3848_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_3856_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3855_wire_constant, tmp_var);
      BITSEL_u8_u1_3856_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_3864_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3863_wire_constant, tmp_var);
      BITSEL_u8_u1_3864_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_3872_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3871_wire_constant, tmp_var);
      BITSEL_u8_u1_3872_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_3880_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3879_wire_constant, tmp_var);
      BITSEL_u8_u1_3880_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_3888_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3887_wire_constant, tmp_var);
      BITSEL_u8_u1_3888_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_3896_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3895_wire_constant, tmp_var);
      BITSEL_u8_u1_3896_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_3904_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3903_wire_constant, tmp_var);
      BITSEL_u8_u1_3904_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_3912_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3911_wire_constant, tmp_var);
      BITSEL_u8_u1_3912_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_3920_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3919_wire_constant, tmp_var);
      BITSEL_u8_u1_3920_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_3928_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3927_wire_constant, tmp_var);
      BITSEL_u8_u1_3928_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_3936_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3935_wire_constant, tmp_var);
      BITSEL_u8_u1_3936_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_3944_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3943_wire_constant, tmp_var);
      BITSEL_u8_u1_3944_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_3952_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3951_wire_constant, tmp_var);
      BITSEL_u8_u1_3952_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_3960_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3959_wire_constant, tmp_var);
      BITSEL_u8_u1_3960_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_3968_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3967_wire_constant, tmp_var);
      BITSEL_u8_u1_3968_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_3976_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3975_wire_constant, tmp_var);
      BITSEL_u8_u1_3976_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_3984_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3983_wire_constant, tmp_var);
      BITSEL_u8_u1_3984_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_3992_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3991_wire_constant, tmp_var);
      BITSEL_u8_u1_3992_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4000_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_3999_wire_constant, tmp_var);
      BITSEL_u8_u1_4000_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4008_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4007_wire_constant, tmp_var);
      BITSEL_u8_u1_4008_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4016_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4015_wire_constant, tmp_var);
      BITSEL_u8_u1_4016_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4024_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4023_wire_constant, tmp_var);
      BITSEL_u8_u1_4024_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4032_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4031_wire_constant, tmp_var);
      BITSEL_u8_u1_4032_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4040_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4039_wire_constant, tmp_var);
      BITSEL_u8_u1_4040_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4048_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4047_wire_constant, tmp_var);
      BITSEL_u8_u1_4048_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4056_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4055_wire_constant, tmp_var);
      BITSEL_u8_u1_4056_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4064_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4063_wire_constant, tmp_var);
      BITSEL_u8_u1_4064_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4072_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4071_wire_constant, tmp_var);
      BITSEL_u8_u1_4072_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4080_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4079_wire_constant, tmp_var);
      BITSEL_u8_u1_4080_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4088_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4087_wire_constant, tmp_var);
      BITSEL_u8_u1_4088_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4096_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4095_wire_constant, tmp_var);
      BITSEL_u8_u1_4096_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4104_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4103_wire_constant, tmp_var);
      BITSEL_u8_u1_4104_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4112_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4111_wire_constant, tmp_var);
      BITSEL_u8_u1_4112_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4120_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4119_wire_constant, tmp_var);
      BITSEL_u8_u1_4120_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4128_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4127_wire_constant, tmp_var);
      BITSEL_u8_u1_4128_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4136_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4135_wire_constant, tmp_var);
      BITSEL_u8_u1_4136_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4144_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4143_wire_constant, tmp_var);
      BITSEL_u8_u1_4144_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4152_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4151_wire_constant, tmp_var);
      BITSEL_u8_u1_4152_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4160_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4159_wire_constant, tmp_var);
      BITSEL_u8_u1_4160_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4168_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4167_wire_constant, tmp_var);
      BITSEL_u8_u1_4168_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4176_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4175_wire_constant, tmp_var);
      BITSEL_u8_u1_4176_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4184_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4183_wire_constant, tmp_var);
      BITSEL_u8_u1_4184_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4192_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4191_wire_constant, tmp_var);
      BITSEL_u8_u1_4192_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4200_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4199_wire_constant, tmp_var);
      BITSEL_u8_u1_4200_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4208_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4207_wire_constant, tmp_var);
      BITSEL_u8_u1_4208_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4216_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4215_wire_constant, tmp_var);
      BITSEL_u8_u1_4216_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4224_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4223_wire_constant, tmp_var);
      BITSEL_u8_u1_4224_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4232_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4231_wire_constant, tmp_var);
      BITSEL_u8_u1_4232_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4240_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4239_wire_constant, tmp_var);
      BITSEL_u8_u1_4240_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4248_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4247_wire_constant, tmp_var);
      BITSEL_u8_u1_4248_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4256_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4255_wire_constant, tmp_var);
      BITSEL_u8_u1_4256_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4264_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4263_wire_constant, tmp_var);
      BITSEL_u8_u1_4264_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4272_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4271_wire_constant, tmp_var);
      BITSEL_u8_u1_4272_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4280_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4279_wire_constant, tmp_var);
      BITSEL_u8_u1_4280_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4288_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4287_wire_constant, tmp_var);
      BITSEL_u8_u1_4288_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4296_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4295_wire_constant, tmp_var);
      BITSEL_u8_u1_4296_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4304_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4303_wire_constant, tmp_var);
      BITSEL_u8_u1_4304_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4312_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4311_wire_constant, tmp_var);
      BITSEL_u8_u1_4312_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4320_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4319_wire_constant, tmp_var);
      BITSEL_u8_u1_4320_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4328_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4327_wire_constant, tmp_var);
      BITSEL_u8_u1_4328_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4336_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4335_wire_constant, tmp_var);
      BITSEL_u8_u1_4336_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4344_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4343_wire_constant, tmp_var);
      BITSEL_u8_u1_4344_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4352_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4351_wire_constant, tmp_var);
      BITSEL_u8_u1_4352_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4360_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4359_wire_constant, tmp_var);
      BITSEL_u8_u1_4360_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4368_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4367_wire_constant, tmp_var);
      BITSEL_u8_u1_4368_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4376_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4375_wire_constant, tmp_var);
      BITSEL_u8_u1_4376_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4384_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4383_wire_constant, tmp_var);
      BITSEL_u8_u1_4384_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4392_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4391_wire_constant, tmp_var);
      BITSEL_u8_u1_4392_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4400_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4399_wire_constant, tmp_var);
      BITSEL_u8_u1_4400_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4408_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4407_wire_constant, tmp_var);
      BITSEL_u8_u1_4408_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4416_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4415_wire_constant, tmp_var);
      BITSEL_u8_u1_4416_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4424_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4423_wire_constant, tmp_var);
      BITSEL_u8_u1_4424_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4432_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4431_wire_constant, tmp_var);
      BITSEL_u8_u1_4432_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4440_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4439_wire_constant, tmp_var);
      BITSEL_u8_u1_4440_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4448_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4447_wire_constant, tmp_var);
      BITSEL_u8_u1_4448_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4456_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4455_wire_constant, tmp_var);
      BITSEL_u8_u1_4456_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4464_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4463_wire_constant, tmp_var);
      BITSEL_u8_u1_4464_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4472_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4471_wire_constant, tmp_var);
      BITSEL_u8_u1_4472_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4480_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4479_wire_constant, tmp_var);
      BITSEL_u8_u1_4480_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4488_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4487_wire_constant, tmp_var);
      BITSEL_u8_u1_4488_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4496_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4495_wire_constant, tmp_var);
      BITSEL_u8_u1_4496_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4504_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4503_wire_constant, tmp_var);
      BITSEL_u8_u1_4504_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4512_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4511_wire_constant, tmp_var);
      BITSEL_u8_u1_4512_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4520_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4519_wire_constant, tmp_var);
      BITSEL_u8_u1_4520_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4528_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4527_wire_constant, tmp_var);
      BITSEL_u8_u1_4528_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4536_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4535_wire_constant, tmp_var);
      BITSEL_u8_u1_4536_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4544_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4543_wire_constant, tmp_var);
      BITSEL_u8_u1_4544_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4552_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4551_wire_constant, tmp_var);
      BITSEL_u8_u1_4552_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4560_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4559_wire_constant, tmp_var);
      BITSEL_u8_u1_4560_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4568_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4567_wire_constant, tmp_var);
      BITSEL_u8_u1_4568_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4576_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4575_wire_constant, tmp_var);
      BITSEL_u8_u1_4576_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4584_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4583_wire_constant, tmp_var);
      BITSEL_u8_u1_4584_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4592_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4591_wire_constant, tmp_var);
      BITSEL_u8_u1_4592_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4600_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4599_wire_constant, tmp_var);
      BITSEL_u8_u1_4600_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4608_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4607_wire_constant, tmp_var);
      BITSEL_u8_u1_4608_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4616_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4615_wire_constant, tmp_var);
      BITSEL_u8_u1_4616_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4624_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4623_wire_constant, tmp_var);
      BITSEL_u8_u1_4624_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4632_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4631_wire_constant, tmp_var);
      BITSEL_u8_u1_4632_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4640_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4639_wire_constant, tmp_var);
      BITSEL_u8_u1_4640_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4648_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4647_wire_constant, tmp_var);
      BITSEL_u8_u1_4648_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4656_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4655_wire_constant, tmp_var);
      BITSEL_u8_u1_4656_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4664_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4663_wire_constant, tmp_var);
      BITSEL_u8_u1_4664_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4672_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4671_wire_constant, tmp_var);
      BITSEL_u8_u1_4672_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4680_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4679_wire_constant, tmp_var);
      BITSEL_u8_u1_4680_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4688_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4687_wire_constant, tmp_var);
      BITSEL_u8_u1_4688_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4696_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4695_wire_constant, tmp_var);
      BITSEL_u8_u1_4696_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4704_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4703_wire_constant, tmp_var);
      BITSEL_u8_u1_4704_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4712_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4711_wire_constant, tmp_var);
      BITSEL_u8_u1_4712_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4720_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4719_wire_constant, tmp_var);
      BITSEL_u8_u1_4720_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4728_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4727_wire_constant, tmp_var);
      BITSEL_u8_u1_4728_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4736_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4735_wire_constant, tmp_var);
      BITSEL_u8_u1_4736_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4744_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4743_wire_constant, tmp_var);
      BITSEL_u8_u1_4744_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4752_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4751_wire_constant, tmp_var);
      BITSEL_u8_u1_4752_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4760_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4759_wire_constant, tmp_var);
      BITSEL_u8_u1_4760_wire <= tmp_var; -- 
    end process;
    -- 
  end Block; -- data_path
  -- 
end Inv_Sbox_2_Volatile_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library work;
use work.ahir_system_global_package.all;
entity Inv_Sbox_3_Volatile is -- 
  port ( -- 
    s_in : in  std_logic_vector(7 downto 0);
    s_out : out  std_logic_vector(7 downto 0)-- 
  );
  -- 
end entity Inv_Sbox_3_Volatile;
architecture Inv_Sbox_3_Volatile_arch of Inv_Sbox_3_Volatile is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector(8-1 downto 0);
  signal default_zero_sig: std_logic;
  -- input port buffer signals
  signal s_in_buffer :  std_logic_vector(7 downto 0);
  -- output port buffer signals
  signal s_out_buffer :  std_logic_vector(7 downto 0);
  -- volatile/operator module components. 
  -- 
begin --  
  -- input handling ------------------------------------------------
  s_in_buffer <= s_in;
  -- output handling  -------------------------------------------------------
  s_out <= s_out_buffer;
  -- the control path --------------------------------------------------
  default_zero_sig <= '0';
  -- volatile module, no control path
  -- the data path
  data_path: Block -- 
    signal BITSEL_u8_u1_4772_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4782_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4792_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4802_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4812_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4822_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4832_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4842_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4852_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4862_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4872_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4882_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4892_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4902_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4912_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4922_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4932_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4942_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4952_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4962_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4972_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4982_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_4992_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5002_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5012_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5022_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5032_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5042_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5052_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5062_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5072_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5082_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5092_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5102_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5112_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5122_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5132_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5142_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5152_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5162_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5172_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5182_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5192_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5202_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5212_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5222_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5232_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5242_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5252_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5262_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5272_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5282_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5292_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5302_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5312_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5322_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5332_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5342_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5352_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5362_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5372_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5382_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5392_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5402_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5412_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5422_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5432_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5442_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5452_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5462_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5472_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5482_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5492_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5502_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5512_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5522_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5532_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5542_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5552_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5562_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5572_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5582_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5592_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5602_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5612_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5622_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5632_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5642_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5652_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5662_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5672_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5682_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5692_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5702_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5712_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5722_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5732_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5742_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5752_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5762_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5772_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5782_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5792_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5802_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5812_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5822_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5832_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5842_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5852_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5862_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5872_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5882_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5892_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5902_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5912_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5922_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5932_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5942_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5952_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5962_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5972_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5982_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_5992_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6002_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6012_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6022_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6032_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6042_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6052_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6060_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6068_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6076_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6084_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6092_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6100_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6108_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6116_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6124_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6132_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6140_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6148_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6156_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6164_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6172_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6180_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6188_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6196_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6204_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6212_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6220_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6228_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6236_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6244_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6252_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6260_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6268_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6276_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6284_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6292_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6300_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6308_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6316_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6324_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6332_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6340_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6348_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6356_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6364_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6372_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6380_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6388_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6396_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6404_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6412_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6420_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6428_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6436_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6444_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6452_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6460_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6468_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6476_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6484_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6492_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6500_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6508_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6516_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6524_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6532_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6540_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6548_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6556_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6564_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6572_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6580_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6588_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6596_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6604_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6612_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6620_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6628_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6636_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6644_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6652_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6660_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6668_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6676_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6684_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6692_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6700_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6708_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6716_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6724_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6732_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6740_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6748_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6756_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6764_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6772_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6780_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6788_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6796_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6804_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6812_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6820_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6828_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6836_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6844_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6852_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6860_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6868_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6876_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6884_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6892_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6900_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6908_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6916_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6924_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6932_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6940_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6948_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6956_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6964_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6972_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6980_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6988_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_6996_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7004_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7012_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7020_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7028_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7036_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7044_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7052_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7060_wire : std_logic_vector(0 downto 0);
    signal IMA0_4778 : std_logic_vector(7 downto 0);
    signal IMA100_5778 : std_logic_vector(7 downto 0);
    signal IMA101_5788 : std_logic_vector(7 downto 0);
    signal IMA102_5798 : std_logic_vector(7 downto 0);
    signal IMA103_5808 : std_logic_vector(7 downto 0);
    signal IMA104_5818 : std_logic_vector(7 downto 0);
    signal IMA105_5828 : std_logic_vector(7 downto 0);
    signal IMA106_5838 : std_logic_vector(7 downto 0);
    signal IMA107_5848 : std_logic_vector(7 downto 0);
    signal IMA108_5858 : std_logic_vector(7 downto 0);
    signal IMA109_5868 : std_logic_vector(7 downto 0);
    signal IMA10_4878 : std_logic_vector(7 downto 0);
    signal IMA110_5878 : std_logic_vector(7 downto 0);
    signal IMA111_5888 : std_logic_vector(7 downto 0);
    signal IMA112_5898 : std_logic_vector(7 downto 0);
    signal IMA113_5908 : std_logic_vector(7 downto 0);
    signal IMA114_5918 : std_logic_vector(7 downto 0);
    signal IMA115_5928 : std_logic_vector(7 downto 0);
    signal IMA116_5938 : std_logic_vector(7 downto 0);
    signal IMA117_5948 : std_logic_vector(7 downto 0);
    signal IMA118_5958 : std_logic_vector(7 downto 0);
    signal IMA119_5968 : std_logic_vector(7 downto 0);
    signal IMA11_4888 : std_logic_vector(7 downto 0);
    signal IMA120_5978 : std_logic_vector(7 downto 0);
    signal IMA121_5988 : std_logic_vector(7 downto 0);
    signal IMA122_5998 : std_logic_vector(7 downto 0);
    signal IMA123_6008 : std_logic_vector(7 downto 0);
    signal IMA124_6018 : std_logic_vector(7 downto 0);
    signal IMA125_6028 : std_logic_vector(7 downto 0);
    signal IMA126_6038 : std_logic_vector(7 downto 0);
    signal IMA127_6048 : std_logic_vector(7 downto 0);
    signal IMA12_4898 : std_logic_vector(7 downto 0);
    signal IMA13_4908 : std_logic_vector(7 downto 0);
    signal IMA14_4918 : std_logic_vector(7 downto 0);
    signal IMA15_4928 : std_logic_vector(7 downto 0);
    signal IMA16_4938 : std_logic_vector(7 downto 0);
    signal IMA17_4948 : std_logic_vector(7 downto 0);
    signal IMA18_4958 : std_logic_vector(7 downto 0);
    signal IMA19_4968 : std_logic_vector(7 downto 0);
    signal IMA1_4788 : std_logic_vector(7 downto 0);
    signal IMA20_4978 : std_logic_vector(7 downto 0);
    signal IMA21_4988 : std_logic_vector(7 downto 0);
    signal IMA22_4998 : std_logic_vector(7 downto 0);
    signal IMA23_5008 : std_logic_vector(7 downto 0);
    signal IMA24_5018 : std_logic_vector(7 downto 0);
    signal IMA25_5028 : std_logic_vector(7 downto 0);
    signal IMA26_5038 : std_logic_vector(7 downto 0);
    signal IMA27_5048 : std_logic_vector(7 downto 0);
    signal IMA28_5058 : std_logic_vector(7 downto 0);
    signal IMA29_5068 : std_logic_vector(7 downto 0);
    signal IMA2_4798 : std_logic_vector(7 downto 0);
    signal IMA30_5078 : std_logic_vector(7 downto 0);
    signal IMA31_5088 : std_logic_vector(7 downto 0);
    signal IMA32_5098 : std_logic_vector(7 downto 0);
    signal IMA33_5108 : std_logic_vector(7 downto 0);
    signal IMA34_5118 : std_logic_vector(7 downto 0);
    signal IMA35_5128 : std_logic_vector(7 downto 0);
    signal IMA36_5138 : std_logic_vector(7 downto 0);
    signal IMA37_5148 : std_logic_vector(7 downto 0);
    signal IMA38_5158 : std_logic_vector(7 downto 0);
    signal IMA39_5168 : std_logic_vector(7 downto 0);
    signal IMA3_4808 : std_logic_vector(7 downto 0);
    signal IMA40_5178 : std_logic_vector(7 downto 0);
    signal IMA41_5188 : std_logic_vector(7 downto 0);
    signal IMA42_5198 : std_logic_vector(7 downto 0);
    signal IMA43_5208 : std_logic_vector(7 downto 0);
    signal IMA44_5218 : std_logic_vector(7 downto 0);
    signal IMA45_5228 : std_logic_vector(7 downto 0);
    signal IMA46_5238 : std_logic_vector(7 downto 0);
    signal IMA47_5248 : std_logic_vector(7 downto 0);
    signal IMA48_5258 : std_logic_vector(7 downto 0);
    signal IMA49_5268 : std_logic_vector(7 downto 0);
    signal IMA4_4818 : std_logic_vector(7 downto 0);
    signal IMA50_5278 : std_logic_vector(7 downto 0);
    signal IMA51_5288 : std_logic_vector(7 downto 0);
    signal IMA52_5298 : std_logic_vector(7 downto 0);
    signal IMA53_5308 : std_logic_vector(7 downto 0);
    signal IMA54_5318 : std_logic_vector(7 downto 0);
    signal IMA55_5328 : std_logic_vector(7 downto 0);
    signal IMA56_5338 : std_logic_vector(7 downto 0);
    signal IMA57_5348 : std_logic_vector(7 downto 0);
    signal IMA58_5358 : std_logic_vector(7 downto 0);
    signal IMA59_5368 : std_logic_vector(7 downto 0);
    signal IMA5_4828 : std_logic_vector(7 downto 0);
    signal IMA60_5378 : std_logic_vector(7 downto 0);
    signal IMA61_5388 : std_logic_vector(7 downto 0);
    signal IMA62_5398 : std_logic_vector(7 downto 0);
    signal IMA63_5408 : std_logic_vector(7 downto 0);
    signal IMA64_5418 : std_logic_vector(7 downto 0);
    signal IMA65_5428 : std_logic_vector(7 downto 0);
    signal IMA66_5438 : std_logic_vector(7 downto 0);
    signal IMA67_5448 : std_logic_vector(7 downto 0);
    signal IMA68_5458 : std_logic_vector(7 downto 0);
    signal IMA69_5468 : std_logic_vector(7 downto 0);
    signal IMA6_4838 : std_logic_vector(7 downto 0);
    signal IMA70_5478 : std_logic_vector(7 downto 0);
    signal IMA71_5488 : std_logic_vector(7 downto 0);
    signal IMA72_5498 : std_logic_vector(7 downto 0);
    signal IMA73_5508 : std_logic_vector(7 downto 0);
    signal IMA74_5518 : std_logic_vector(7 downto 0);
    signal IMA75_5528 : std_logic_vector(7 downto 0);
    signal IMA76_5538 : std_logic_vector(7 downto 0);
    signal IMA77_5548 : std_logic_vector(7 downto 0);
    signal IMA78_5558 : std_logic_vector(7 downto 0);
    signal IMA79_5568 : std_logic_vector(7 downto 0);
    signal IMA7_4848 : std_logic_vector(7 downto 0);
    signal IMA80_5578 : std_logic_vector(7 downto 0);
    signal IMA81_5588 : std_logic_vector(7 downto 0);
    signal IMA82_5598 : std_logic_vector(7 downto 0);
    signal IMA83_5608 : std_logic_vector(7 downto 0);
    signal IMA84_5618 : std_logic_vector(7 downto 0);
    signal IMA85_5628 : std_logic_vector(7 downto 0);
    signal IMA86_5638 : std_logic_vector(7 downto 0);
    signal IMA87_5648 : std_logic_vector(7 downto 0);
    signal IMA88_5658 : std_logic_vector(7 downto 0);
    signal IMA89_5668 : std_logic_vector(7 downto 0);
    signal IMA8_4858 : std_logic_vector(7 downto 0);
    signal IMA90_5678 : std_logic_vector(7 downto 0);
    signal IMA91_5688 : std_logic_vector(7 downto 0);
    signal IMA92_5698 : std_logic_vector(7 downto 0);
    signal IMA93_5708 : std_logic_vector(7 downto 0);
    signal IMA94_5718 : std_logic_vector(7 downto 0);
    signal IMA95_5728 : std_logic_vector(7 downto 0);
    signal IMA96_5738 : std_logic_vector(7 downto 0);
    signal IMA97_5748 : std_logic_vector(7 downto 0);
    signal IMA98_5758 : std_logic_vector(7 downto 0);
    signal IMA99_5768 : std_logic_vector(7 downto 0);
    signal IMA9_4868 : std_logic_vector(7 downto 0);
    signal IMB0_6056 : std_logic_vector(7 downto 0);
    signal IMB10_6136 : std_logic_vector(7 downto 0);
    signal IMB11_6144 : std_logic_vector(7 downto 0);
    signal IMB12_6152 : std_logic_vector(7 downto 0);
    signal IMB13_6160 : std_logic_vector(7 downto 0);
    signal IMB14_6168 : std_logic_vector(7 downto 0);
    signal IMB15_6176 : std_logic_vector(7 downto 0);
    signal IMB16_6184 : std_logic_vector(7 downto 0);
    signal IMB17_6192 : std_logic_vector(7 downto 0);
    signal IMB18_6200 : std_logic_vector(7 downto 0);
    signal IMB19_6208 : std_logic_vector(7 downto 0);
    signal IMB1_6064 : std_logic_vector(7 downto 0);
    signal IMB20_6216 : std_logic_vector(7 downto 0);
    signal IMB21_6224 : std_logic_vector(7 downto 0);
    signal IMB22_6232 : std_logic_vector(7 downto 0);
    signal IMB23_6240 : std_logic_vector(7 downto 0);
    signal IMB24_6248 : std_logic_vector(7 downto 0);
    signal IMB25_6256 : std_logic_vector(7 downto 0);
    signal IMB26_6264 : std_logic_vector(7 downto 0);
    signal IMB27_6272 : std_logic_vector(7 downto 0);
    signal IMB28_6280 : std_logic_vector(7 downto 0);
    signal IMB29_6288 : std_logic_vector(7 downto 0);
    signal IMB2_6072 : std_logic_vector(7 downto 0);
    signal IMB30_6296 : std_logic_vector(7 downto 0);
    signal IMB31_6304 : std_logic_vector(7 downto 0);
    signal IMB32_6312 : std_logic_vector(7 downto 0);
    signal IMB33_6320 : std_logic_vector(7 downto 0);
    signal IMB34_6328 : std_logic_vector(7 downto 0);
    signal IMB35_6336 : std_logic_vector(7 downto 0);
    signal IMB36_6344 : std_logic_vector(7 downto 0);
    signal IMB37_6352 : std_logic_vector(7 downto 0);
    signal IMB38_6360 : std_logic_vector(7 downto 0);
    signal IMB39_6368 : std_logic_vector(7 downto 0);
    signal IMB3_6080 : std_logic_vector(7 downto 0);
    signal IMB40_6376 : std_logic_vector(7 downto 0);
    signal IMB41_6384 : std_logic_vector(7 downto 0);
    signal IMB42_6392 : std_logic_vector(7 downto 0);
    signal IMB43_6400 : std_logic_vector(7 downto 0);
    signal IMB44_6408 : std_logic_vector(7 downto 0);
    signal IMB45_6416 : std_logic_vector(7 downto 0);
    signal IMB46_6424 : std_logic_vector(7 downto 0);
    signal IMB47_6432 : std_logic_vector(7 downto 0);
    signal IMB48_6440 : std_logic_vector(7 downto 0);
    signal IMB49_6448 : std_logic_vector(7 downto 0);
    signal IMB4_6088 : std_logic_vector(7 downto 0);
    signal IMB50_6456 : std_logic_vector(7 downto 0);
    signal IMB51_6464 : std_logic_vector(7 downto 0);
    signal IMB52_6472 : std_logic_vector(7 downto 0);
    signal IMB53_6480 : std_logic_vector(7 downto 0);
    signal IMB54_6488 : std_logic_vector(7 downto 0);
    signal IMB55_6496 : std_logic_vector(7 downto 0);
    signal IMB56_6504 : std_logic_vector(7 downto 0);
    signal IMB57_6512 : std_logic_vector(7 downto 0);
    signal IMB58_6520 : std_logic_vector(7 downto 0);
    signal IMB59_6528 : std_logic_vector(7 downto 0);
    signal IMB5_6096 : std_logic_vector(7 downto 0);
    signal IMB60_6536 : std_logic_vector(7 downto 0);
    signal IMB61_6544 : std_logic_vector(7 downto 0);
    signal IMB62_6552 : std_logic_vector(7 downto 0);
    signal IMB63_6560 : std_logic_vector(7 downto 0);
    signal IMB6_6104 : std_logic_vector(7 downto 0);
    signal IMB7_6112 : std_logic_vector(7 downto 0);
    signal IMB8_6120 : std_logic_vector(7 downto 0);
    signal IMB9_6128 : std_logic_vector(7 downto 0);
    signal IMC0_6568 : std_logic_vector(7 downto 0);
    signal IMC10_6648 : std_logic_vector(7 downto 0);
    signal IMC11_6656 : std_logic_vector(7 downto 0);
    signal IMC12_6664 : std_logic_vector(7 downto 0);
    signal IMC13_6672 : std_logic_vector(7 downto 0);
    signal IMC14_6680 : std_logic_vector(7 downto 0);
    signal IMC15_6688 : std_logic_vector(7 downto 0);
    signal IMC16_6696 : std_logic_vector(7 downto 0);
    signal IMC17_6704 : std_logic_vector(7 downto 0);
    signal IMC18_6712 : std_logic_vector(7 downto 0);
    signal IMC19_6720 : std_logic_vector(7 downto 0);
    signal IMC1_6576 : std_logic_vector(7 downto 0);
    signal IMC20_6728 : std_logic_vector(7 downto 0);
    signal IMC21_6736 : std_logic_vector(7 downto 0);
    signal IMC22_6744 : std_logic_vector(7 downto 0);
    signal IMC23_6752 : std_logic_vector(7 downto 0);
    signal IMC24_6760 : std_logic_vector(7 downto 0);
    signal IMC25_6768 : std_logic_vector(7 downto 0);
    signal IMC26_6776 : std_logic_vector(7 downto 0);
    signal IMC27_6784 : std_logic_vector(7 downto 0);
    signal IMC28_6792 : std_logic_vector(7 downto 0);
    signal IMC29_6800 : std_logic_vector(7 downto 0);
    signal IMC2_6584 : std_logic_vector(7 downto 0);
    signal IMC30_6808 : std_logic_vector(7 downto 0);
    signal IMC31_6816 : std_logic_vector(7 downto 0);
    signal IMC3_6592 : std_logic_vector(7 downto 0);
    signal IMC4_6600 : std_logic_vector(7 downto 0);
    signal IMC5_6608 : std_logic_vector(7 downto 0);
    signal IMC6_6616 : std_logic_vector(7 downto 0);
    signal IMC7_6624 : std_logic_vector(7 downto 0);
    signal IMC8_6632 : std_logic_vector(7 downto 0);
    signal IMC9_6640 : std_logic_vector(7 downto 0);
    signal IMD0_6824 : std_logic_vector(7 downto 0);
    signal IMD10_6904 : std_logic_vector(7 downto 0);
    signal IMD11_6912 : std_logic_vector(7 downto 0);
    signal IMD12_6920 : std_logic_vector(7 downto 0);
    signal IMD13_6928 : std_logic_vector(7 downto 0);
    signal IMD14_6936 : std_logic_vector(7 downto 0);
    signal IMD15_6944 : std_logic_vector(7 downto 0);
    signal IMD1_6832 : std_logic_vector(7 downto 0);
    signal IMD2_6840 : std_logic_vector(7 downto 0);
    signal IMD3_6848 : std_logic_vector(7 downto 0);
    signal IMD4_6856 : std_logic_vector(7 downto 0);
    signal IMD5_6864 : std_logic_vector(7 downto 0);
    signal IMD6_6872 : std_logic_vector(7 downto 0);
    signal IMD7_6880 : std_logic_vector(7 downto 0);
    signal IMD8_6888 : std_logic_vector(7 downto 0);
    signal IMD9_6896 : std_logic_vector(7 downto 0);
    signal IME0_6952 : std_logic_vector(7 downto 0);
    signal IME1_6960 : std_logic_vector(7 downto 0);
    signal IME2_6968 : std_logic_vector(7 downto 0);
    signal IME3_6976 : std_logic_vector(7 downto 0);
    signal IME4_6984 : std_logic_vector(7 downto 0);
    signal IME5_6992 : std_logic_vector(7 downto 0);
    signal IME6_7000 : std_logic_vector(7 downto 0);
    signal IME7_7008 : std_logic_vector(7 downto 0);
    signal IMF0_7016 : std_logic_vector(7 downto 0);
    signal IMF1_7024 : std_logic_vector(7 downto 0);
    signal IMF2_7032 : std_logic_vector(7 downto 0);
    signal IMF3_7040 : std_logic_vector(7 downto 0);
    signal IMG0_7048 : std_logic_vector(7 downto 0);
    signal IMG1_7056 : std_logic_vector(7 downto 0);
    signal konst_4771_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4781_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4791_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4801_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4811_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4821_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4831_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4841_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4851_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4861_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4871_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4881_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4891_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4901_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4911_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4921_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4931_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4941_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4951_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4961_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4971_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4981_wire_constant : std_logic_vector(7 downto 0);
    signal konst_4991_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5001_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5011_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5021_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5031_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5041_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5051_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5061_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5071_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5081_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5091_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5101_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5111_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5121_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5131_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5141_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5151_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5161_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5171_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5181_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5191_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5201_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5211_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5221_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5231_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5241_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5251_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5261_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5271_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5281_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5291_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5301_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5311_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5321_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5331_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5341_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5351_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5361_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5371_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5381_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5391_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5401_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5411_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5421_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5431_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5441_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5451_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5461_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5471_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5481_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5491_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5501_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5511_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5521_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5531_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5541_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5551_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5561_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5571_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5581_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5591_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5601_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5611_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5621_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5631_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5641_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5651_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5661_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5671_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5681_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5691_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5701_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5711_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5721_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5731_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5741_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5751_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5761_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5771_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5781_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5791_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5801_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5811_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5821_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5831_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5841_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5851_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5861_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5871_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5881_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5891_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5901_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5911_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5921_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5931_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5941_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5951_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5961_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5971_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5981_wire_constant : std_logic_vector(7 downto 0);
    signal konst_5991_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6001_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6011_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6021_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6031_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6041_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6051_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6059_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6067_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6075_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6083_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6091_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6099_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6107_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6115_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6123_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6131_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6139_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6147_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6155_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6163_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6171_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6179_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6187_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6195_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6203_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6211_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6219_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6227_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6235_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6243_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6251_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6259_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6267_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6275_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6283_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6291_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6299_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6307_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6315_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6323_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6331_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6339_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6347_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6355_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6363_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6371_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6379_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6387_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6395_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6403_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6411_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6419_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6427_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6435_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6443_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6451_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6459_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6467_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6475_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6483_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6491_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6499_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6507_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6515_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6523_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6531_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6539_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6547_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6555_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6563_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6571_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6579_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6587_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6595_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6603_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6611_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6619_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6627_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6635_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6643_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6651_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6659_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6667_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6675_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6683_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6691_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6699_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6707_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6715_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6723_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6731_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6739_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6747_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6755_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6763_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6771_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6779_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6787_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6795_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6803_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6811_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6819_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6827_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6835_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6843_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6851_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6859_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6867_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6875_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6883_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6891_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6899_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6907_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6915_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6923_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6931_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6939_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6947_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6955_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6963_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6971_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6979_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6987_wire_constant : std_logic_vector(7 downto 0);
    signal konst_6995_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7003_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7011_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7019_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7027_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7035_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7043_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7051_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7059_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4774_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4776_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4784_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4786_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4794_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4796_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4804_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4806_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4814_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4816_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4824_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4826_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4834_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4836_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4844_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4846_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4854_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4856_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4864_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4866_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4874_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4876_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4884_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4886_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4894_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4896_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4904_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4906_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4914_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4916_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4924_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4926_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4934_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4936_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4944_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4946_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4954_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4956_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4964_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4966_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4974_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4976_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4984_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4986_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4994_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_4996_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5004_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5006_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5014_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5016_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5024_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5026_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5034_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5036_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5044_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5046_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5054_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5056_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5064_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5066_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5074_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5076_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5084_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5086_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5094_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5096_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5104_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5106_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5114_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5116_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5124_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5126_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5134_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5136_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5144_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5146_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5154_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5156_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5164_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5166_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5174_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5176_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5184_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5186_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5194_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5196_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5204_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5206_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5214_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5216_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5224_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5226_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5234_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5236_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5244_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5246_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5254_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5256_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5264_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5266_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5274_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5276_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5284_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5286_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5294_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5296_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5304_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5306_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5314_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5316_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5324_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5326_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5334_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5336_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5344_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5346_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5354_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5356_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5364_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5366_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5374_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5376_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5384_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5386_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5394_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5396_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5404_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5406_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5414_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5416_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5424_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5426_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5434_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5436_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5444_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5446_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5454_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5456_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5464_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5466_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5474_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5476_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5484_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5486_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5494_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5496_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5504_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5506_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5514_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5516_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5524_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5526_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5534_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5536_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5544_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5546_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5554_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5556_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5564_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5566_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5574_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5576_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5584_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5586_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5594_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5596_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5604_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5606_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5614_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5616_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5624_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5626_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5634_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5636_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5644_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5646_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5654_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5656_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5664_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5666_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5674_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5676_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5684_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5686_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5694_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5696_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5704_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5706_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5714_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5716_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5724_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5726_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5734_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5736_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5744_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5746_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5754_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5756_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5764_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5766_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5774_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5776_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5784_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5786_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5794_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5796_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5804_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5806_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5814_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5816_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5824_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5826_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5834_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5836_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5844_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5846_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5854_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5856_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5864_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5866_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5874_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5876_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5884_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5886_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5894_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5896_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5904_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5906_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5914_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5916_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5924_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5926_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5934_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5936_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5944_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5946_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5954_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5956_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5964_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5966_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5974_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5976_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5984_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5986_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5994_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_5996_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_6004_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_6006_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_6014_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_6016_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_6024_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_6026_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_6034_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_6036_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_6044_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_6046_wire_constant : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    konst_4771_wire_constant <= "00000000";
    konst_4781_wire_constant <= "00000000";
    konst_4791_wire_constant <= "00000000";
    konst_4801_wire_constant <= "00000000";
    konst_4811_wire_constant <= "00000000";
    konst_4821_wire_constant <= "00000000";
    konst_4831_wire_constant <= "00000000";
    konst_4841_wire_constant <= "00000000";
    konst_4851_wire_constant <= "00000000";
    konst_4861_wire_constant <= "00000000";
    konst_4871_wire_constant <= "00000000";
    konst_4881_wire_constant <= "00000000";
    konst_4891_wire_constant <= "00000000";
    konst_4901_wire_constant <= "00000000";
    konst_4911_wire_constant <= "00000000";
    konst_4921_wire_constant <= "00000000";
    konst_4931_wire_constant <= "00000000";
    konst_4941_wire_constant <= "00000000";
    konst_4951_wire_constant <= "00000000";
    konst_4961_wire_constant <= "00000000";
    konst_4971_wire_constant <= "00000000";
    konst_4981_wire_constant <= "00000000";
    konst_4991_wire_constant <= "00000000";
    konst_5001_wire_constant <= "00000000";
    konst_5011_wire_constant <= "00000000";
    konst_5021_wire_constant <= "00000000";
    konst_5031_wire_constant <= "00000000";
    konst_5041_wire_constant <= "00000000";
    konst_5051_wire_constant <= "00000000";
    konst_5061_wire_constant <= "00000000";
    konst_5071_wire_constant <= "00000000";
    konst_5081_wire_constant <= "00000000";
    konst_5091_wire_constant <= "00000000";
    konst_5101_wire_constant <= "00000000";
    konst_5111_wire_constant <= "00000000";
    konst_5121_wire_constant <= "00000000";
    konst_5131_wire_constant <= "00000000";
    konst_5141_wire_constant <= "00000000";
    konst_5151_wire_constant <= "00000000";
    konst_5161_wire_constant <= "00000000";
    konst_5171_wire_constant <= "00000000";
    konst_5181_wire_constant <= "00000000";
    konst_5191_wire_constant <= "00000000";
    konst_5201_wire_constant <= "00000000";
    konst_5211_wire_constant <= "00000000";
    konst_5221_wire_constant <= "00000000";
    konst_5231_wire_constant <= "00000000";
    konst_5241_wire_constant <= "00000000";
    konst_5251_wire_constant <= "00000000";
    konst_5261_wire_constant <= "00000000";
    konst_5271_wire_constant <= "00000000";
    konst_5281_wire_constant <= "00000000";
    konst_5291_wire_constant <= "00000000";
    konst_5301_wire_constant <= "00000000";
    konst_5311_wire_constant <= "00000000";
    konst_5321_wire_constant <= "00000000";
    konst_5331_wire_constant <= "00000000";
    konst_5341_wire_constant <= "00000000";
    konst_5351_wire_constant <= "00000000";
    konst_5361_wire_constant <= "00000000";
    konst_5371_wire_constant <= "00000000";
    konst_5381_wire_constant <= "00000000";
    konst_5391_wire_constant <= "00000000";
    konst_5401_wire_constant <= "00000000";
    konst_5411_wire_constant <= "00000000";
    konst_5421_wire_constant <= "00000000";
    konst_5431_wire_constant <= "00000000";
    konst_5441_wire_constant <= "00000000";
    konst_5451_wire_constant <= "00000000";
    konst_5461_wire_constant <= "00000000";
    konst_5471_wire_constant <= "00000000";
    konst_5481_wire_constant <= "00000000";
    konst_5491_wire_constant <= "00000000";
    konst_5501_wire_constant <= "00000000";
    konst_5511_wire_constant <= "00000000";
    konst_5521_wire_constant <= "00000000";
    konst_5531_wire_constant <= "00000000";
    konst_5541_wire_constant <= "00000000";
    konst_5551_wire_constant <= "00000000";
    konst_5561_wire_constant <= "00000000";
    konst_5571_wire_constant <= "00000000";
    konst_5581_wire_constant <= "00000000";
    konst_5591_wire_constant <= "00000000";
    konst_5601_wire_constant <= "00000000";
    konst_5611_wire_constant <= "00000000";
    konst_5621_wire_constant <= "00000000";
    konst_5631_wire_constant <= "00000000";
    konst_5641_wire_constant <= "00000000";
    konst_5651_wire_constant <= "00000000";
    konst_5661_wire_constant <= "00000000";
    konst_5671_wire_constant <= "00000000";
    konst_5681_wire_constant <= "00000000";
    konst_5691_wire_constant <= "00000000";
    konst_5701_wire_constant <= "00000000";
    konst_5711_wire_constant <= "00000000";
    konst_5721_wire_constant <= "00000000";
    konst_5731_wire_constant <= "00000000";
    konst_5741_wire_constant <= "00000000";
    konst_5751_wire_constant <= "00000000";
    konst_5761_wire_constant <= "00000000";
    konst_5771_wire_constant <= "00000000";
    konst_5781_wire_constant <= "00000000";
    konst_5791_wire_constant <= "00000000";
    konst_5801_wire_constant <= "00000000";
    konst_5811_wire_constant <= "00000000";
    konst_5821_wire_constant <= "00000000";
    konst_5831_wire_constant <= "00000000";
    konst_5841_wire_constant <= "00000000";
    konst_5851_wire_constant <= "00000000";
    konst_5861_wire_constant <= "00000000";
    konst_5871_wire_constant <= "00000000";
    konst_5881_wire_constant <= "00000000";
    konst_5891_wire_constant <= "00000000";
    konst_5901_wire_constant <= "00000000";
    konst_5911_wire_constant <= "00000000";
    konst_5921_wire_constant <= "00000000";
    konst_5931_wire_constant <= "00000000";
    konst_5941_wire_constant <= "00000000";
    konst_5951_wire_constant <= "00000000";
    konst_5961_wire_constant <= "00000000";
    konst_5971_wire_constant <= "00000000";
    konst_5981_wire_constant <= "00000000";
    konst_5991_wire_constant <= "00000000";
    konst_6001_wire_constant <= "00000000";
    konst_6011_wire_constant <= "00000000";
    konst_6021_wire_constant <= "00000000";
    konst_6031_wire_constant <= "00000000";
    konst_6041_wire_constant <= "00000000";
    konst_6051_wire_constant <= "00000001";
    konst_6059_wire_constant <= "00000001";
    konst_6067_wire_constant <= "00000001";
    konst_6075_wire_constant <= "00000001";
    konst_6083_wire_constant <= "00000001";
    konst_6091_wire_constant <= "00000001";
    konst_6099_wire_constant <= "00000001";
    konst_6107_wire_constant <= "00000001";
    konst_6115_wire_constant <= "00000001";
    konst_6123_wire_constant <= "00000001";
    konst_6131_wire_constant <= "00000001";
    konst_6139_wire_constant <= "00000001";
    konst_6147_wire_constant <= "00000001";
    konst_6155_wire_constant <= "00000001";
    konst_6163_wire_constant <= "00000001";
    konst_6171_wire_constant <= "00000001";
    konst_6179_wire_constant <= "00000001";
    konst_6187_wire_constant <= "00000001";
    konst_6195_wire_constant <= "00000001";
    konst_6203_wire_constant <= "00000001";
    konst_6211_wire_constant <= "00000001";
    konst_6219_wire_constant <= "00000001";
    konst_6227_wire_constant <= "00000001";
    konst_6235_wire_constant <= "00000001";
    konst_6243_wire_constant <= "00000001";
    konst_6251_wire_constant <= "00000001";
    konst_6259_wire_constant <= "00000001";
    konst_6267_wire_constant <= "00000001";
    konst_6275_wire_constant <= "00000001";
    konst_6283_wire_constant <= "00000001";
    konst_6291_wire_constant <= "00000001";
    konst_6299_wire_constant <= "00000001";
    konst_6307_wire_constant <= "00000001";
    konst_6315_wire_constant <= "00000001";
    konst_6323_wire_constant <= "00000001";
    konst_6331_wire_constant <= "00000001";
    konst_6339_wire_constant <= "00000001";
    konst_6347_wire_constant <= "00000001";
    konst_6355_wire_constant <= "00000001";
    konst_6363_wire_constant <= "00000001";
    konst_6371_wire_constant <= "00000001";
    konst_6379_wire_constant <= "00000001";
    konst_6387_wire_constant <= "00000001";
    konst_6395_wire_constant <= "00000001";
    konst_6403_wire_constant <= "00000001";
    konst_6411_wire_constant <= "00000001";
    konst_6419_wire_constant <= "00000001";
    konst_6427_wire_constant <= "00000001";
    konst_6435_wire_constant <= "00000001";
    konst_6443_wire_constant <= "00000001";
    konst_6451_wire_constant <= "00000001";
    konst_6459_wire_constant <= "00000001";
    konst_6467_wire_constant <= "00000001";
    konst_6475_wire_constant <= "00000001";
    konst_6483_wire_constant <= "00000001";
    konst_6491_wire_constant <= "00000001";
    konst_6499_wire_constant <= "00000001";
    konst_6507_wire_constant <= "00000001";
    konst_6515_wire_constant <= "00000001";
    konst_6523_wire_constant <= "00000001";
    konst_6531_wire_constant <= "00000001";
    konst_6539_wire_constant <= "00000001";
    konst_6547_wire_constant <= "00000001";
    konst_6555_wire_constant <= "00000001";
    konst_6563_wire_constant <= "00000010";
    konst_6571_wire_constant <= "00000010";
    konst_6579_wire_constant <= "00000010";
    konst_6587_wire_constant <= "00000010";
    konst_6595_wire_constant <= "00000010";
    konst_6603_wire_constant <= "00000010";
    konst_6611_wire_constant <= "00000010";
    konst_6619_wire_constant <= "00000010";
    konst_6627_wire_constant <= "00000010";
    konst_6635_wire_constant <= "00000010";
    konst_6643_wire_constant <= "00000010";
    konst_6651_wire_constant <= "00000010";
    konst_6659_wire_constant <= "00000010";
    konst_6667_wire_constant <= "00000010";
    konst_6675_wire_constant <= "00000010";
    konst_6683_wire_constant <= "00000010";
    konst_6691_wire_constant <= "00000010";
    konst_6699_wire_constant <= "00000010";
    konst_6707_wire_constant <= "00000010";
    konst_6715_wire_constant <= "00000010";
    konst_6723_wire_constant <= "00000010";
    konst_6731_wire_constant <= "00000010";
    konst_6739_wire_constant <= "00000010";
    konst_6747_wire_constant <= "00000010";
    konst_6755_wire_constant <= "00000010";
    konst_6763_wire_constant <= "00000010";
    konst_6771_wire_constant <= "00000010";
    konst_6779_wire_constant <= "00000010";
    konst_6787_wire_constant <= "00000010";
    konst_6795_wire_constant <= "00000010";
    konst_6803_wire_constant <= "00000010";
    konst_6811_wire_constant <= "00000010";
    konst_6819_wire_constant <= "00000011";
    konst_6827_wire_constant <= "00000011";
    konst_6835_wire_constant <= "00000011";
    konst_6843_wire_constant <= "00000011";
    konst_6851_wire_constant <= "00000011";
    konst_6859_wire_constant <= "00000011";
    konst_6867_wire_constant <= "00000011";
    konst_6875_wire_constant <= "00000011";
    konst_6883_wire_constant <= "00000011";
    konst_6891_wire_constant <= "00000011";
    konst_6899_wire_constant <= "00000011";
    konst_6907_wire_constant <= "00000011";
    konst_6915_wire_constant <= "00000011";
    konst_6923_wire_constant <= "00000011";
    konst_6931_wire_constant <= "00000011";
    konst_6939_wire_constant <= "00000011";
    konst_6947_wire_constant <= "00000100";
    konst_6955_wire_constant <= "00000100";
    konst_6963_wire_constant <= "00000100";
    konst_6971_wire_constant <= "00000100";
    konst_6979_wire_constant <= "00000100";
    konst_6987_wire_constant <= "00000100";
    konst_6995_wire_constant <= "00000100";
    konst_7003_wire_constant <= "00000100";
    konst_7011_wire_constant <= "00000101";
    konst_7019_wire_constant <= "00000101";
    konst_7027_wire_constant <= "00000101";
    konst_7035_wire_constant <= "00000101";
    konst_7043_wire_constant <= "00000110";
    konst_7051_wire_constant <= "00000110";
    konst_7059_wire_constant <= "00000111";
    type_cast_4774_wire_constant <= "00001001";
    type_cast_4776_wire_constant <= "01010010";
    type_cast_4784_wire_constant <= "11010101";
    type_cast_4786_wire_constant <= "01101010";
    type_cast_4794_wire_constant <= "00110110";
    type_cast_4796_wire_constant <= "00110000";
    type_cast_4804_wire_constant <= "00111000";
    type_cast_4806_wire_constant <= "10100101";
    type_cast_4814_wire_constant <= "01000000";
    type_cast_4816_wire_constant <= "10111111";
    type_cast_4824_wire_constant <= "10011110";
    type_cast_4826_wire_constant <= "10100011";
    type_cast_4834_wire_constant <= "11110011";
    type_cast_4836_wire_constant <= "10000001";
    type_cast_4844_wire_constant <= "11111011";
    type_cast_4846_wire_constant <= "11010111";
    type_cast_4854_wire_constant <= "11100011";
    type_cast_4856_wire_constant <= "01111100";
    type_cast_4864_wire_constant <= "10000010";
    type_cast_4866_wire_constant <= "00111001";
    type_cast_4874_wire_constant <= "00101111";
    type_cast_4876_wire_constant <= "10011011";
    type_cast_4884_wire_constant <= "10000111";
    type_cast_4886_wire_constant <= "11111111";
    type_cast_4894_wire_constant <= "10001110";
    type_cast_4896_wire_constant <= "00110100";
    type_cast_4904_wire_constant <= "01000100";
    type_cast_4906_wire_constant <= "01000011";
    type_cast_4914_wire_constant <= "11011110";
    type_cast_4916_wire_constant <= "11000100";
    type_cast_4924_wire_constant <= "11001011";
    type_cast_4926_wire_constant <= "11101001";
    type_cast_4934_wire_constant <= "01111011";
    type_cast_4936_wire_constant <= "01010100";
    type_cast_4944_wire_constant <= "00110010";
    type_cast_4946_wire_constant <= "10010100";
    type_cast_4954_wire_constant <= "11000010";
    type_cast_4956_wire_constant <= "10100110";
    type_cast_4964_wire_constant <= "00111101";
    type_cast_4966_wire_constant <= "00100011";
    type_cast_4974_wire_constant <= "01001100";
    type_cast_4976_wire_constant <= "11101110";
    type_cast_4984_wire_constant <= "00001011";
    type_cast_4986_wire_constant <= "10010101";
    type_cast_4994_wire_constant <= "11111010";
    type_cast_4996_wire_constant <= "01000010";
    type_cast_5004_wire_constant <= "01001110";
    type_cast_5006_wire_constant <= "11000011";
    type_cast_5014_wire_constant <= "00101110";
    type_cast_5016_wire_constant <= "00001000";
    type_cast_5024_wire_constant <= "01100110";
    type_cast_5026_wire_constant <= "10100001";
    type_cast_5034_wire_constant <= "11011001";
    type_cast_5036_wire_constant <= "00101000";
    type_cast_5044_wire_constant <= "10110010";
    type_cast_5046_wire_constant <= "00100100";
    type_cast_5054_wire_constant <= "01011011";
    type_cast_5056_wire_constant <= "01110110";
    type_cast_5064_wire_constant <= "01001001";
    type_cast_5066_wire_constant <= "10100010";
    type_cast_5074_wire_constant <= "10001011";
    type_cast_5076_wire_constant <= "01101101";
    type_cast_5084_wire_constant <= "00100101";
    type_cast_5086_wire_constant <= "11010001";
    type_cast_5094_wire_constant <= "11111000";
    type_cast_5096_wire_constant <= "01110010";
    type_cast_5104_wire_constant <= "01100100";
    type_cast_5106_wire_constant <= "11110110";
    type_cast_5114_wire_constant <= "01101000";
    type_cast_5116_wire_constant <= "10000110";
    type_cast_5124_wire_constant <= "00010110";
    type_cast_5126_wire_constant <= "10011000";
    type_cast_5134_wire_constant <= "10100100";
    type_cast_5136_wire_constant <= "11010100";
    type_cast_5144_wire_constant <= "11001100";
    type_cast_5146_wire_constant <= "01011100";
    type_cast_5154_wire_constant <= "01100101";
    type_cast_5156_wire_constant <= "01011101";
    type_cast_5164_wire_constant <= "10010010";
    type_cast_5166_wire_constant <= "10110110";
    type_cast_5174_wire_constant <= "01110000";
    type_cast_5176_wire_constant <= "01101100";
    type_cast_5184_wire_constant <= "01010000";
    type_cast_5186_wire_constant <= "01001000";
    type_cast_5194_wire_constant <= "11101101";
    type_cast_5196_wire_constant <= "11111101";
    type_cast_5204_wire_constant <= "11011010";
    type_cast_5206_wire_constant <= "10111001";
    type_cast_5214_wire_constant <= "00010101";
    type_cast_5216_wire_constant <= "01011110";
    type_cast_5224_wire_constant <= "01010111";
    type_cast_5226_wire_constant <= "01000110";
    type_cast_5234_wire_constant <= "10001101";
    type_cast_5236_wire_constant <= "10100111";
    type_cast_5244_wire_constant <= "10000100";
    type_cast_5246_wire_constant <= "10011101";
    type_cast_5254_wire_constant <= "11011000";
    type_cast_5256_wire_constant <= "10010000";
    type_cast_5264_wire_constant <= "00000000";
    type_cast_5266_wire_constant <= "10101011";
    type_cast_5274_wire_constant <= "10111100";
    type_cast_5276_wire_constant <= "10001100";
    type_cast_5284_wire_constant <= "00001010";
    type_cast_5286_wire_constant <= "11010011";
    type_cast_5294_wire_constant <= "11100100";
    type_cast_5296_wire_constant <= "11110111";
    type_cast_5304_wire_constant <= "00000101";
    type_cast_5306_wire_constant <= "01011000";
    type_cast_5314_wire_constant <= "10110011";
    type_cast_5316_wire_constant <= "10111000";
    type_cast_5324_wire_constant <= "00000110";
    type_cast_5326_wire_constant <= "01000101";
    type_cast_5334_wire_constant <= "00101100";
    type_cast_5336_wire_constant <= "11010000";
    type_cast_5344_wire_constant <= "10001111";
    type_cast_5346_wire_constant <= "00011110";
    type_cast_5354_wire_constant <= "00111111";
    type_cast_5356_wire_constant <= "11001010";
    type_cast_5364_wire_constant <= "00000010";
    type_cast_5366_wire_constant <= "00001111";
    type_cast_5374_wire_constant <= "10101111";
    type_cast_5376_wire_constant <= "11000001";
    type_cast_5384_wire_constant <= "00000011";
    type_cast_5386_wire_constant <= "10111101";
    type_cast_5394_wire_constant <= "00010011";
    type_cast_5396_wire_constant <= "00000001";
    type_cast_5404_wire_constant <= "01101011";
    type_cast_5406_wire_constant <= "10001010";
    type_cast_5414_wire_constant <= "10010001";
    type_cast_5416_wire_constant <= "00111010";
    type_cast_5424_wire_constant <= "01000001";
    type_cast_5426_wire_constant <= "00010001";
    type_cast_5434_wire_constant <= "01100111";
    type_cast_5436_wire_constant <= "01001111";
    type_cast_5444_wire_constant <= "11101010";
    type_cast_5446_wire_constant <= "11011100";
    type_cast_5454_wire_constant <= "11110010";
    type_cast_5456_wire_constant <= "10010111";
    type_cast_5464_wire_constant <= "11001110";
    type_cast_5466_wire_constant <= "11001111";
    type_cast_5474_wire_constant <= "10110100";
    type_cast_5476_wire_constant <= "11110000";
    type_cast_5484_wire_constant <= "01110011";
    type_cast_5486_wire_constant <= "11100110";
    type_cast_5494_wire_constant <= "10101100";
    type_cast_5496_wire_constant <= "10010110";
    type_cast_5504_wire_constant <= "00100010";
    type_cast_5506_wire_constant <= "01110100";
    type_cast_5514_wire_constant <= "10101101";
    type_cast_5516_wire_constant <= "11100111";
    type_cast_5524_wire_constant <= "10000101";
    type_cast_5526_wire_constant <= "00110101";
    type_cast_5534_wire_constant <= "11111001";
    type_cast_5536_wire_constant <= "11100010";
    type_cast_5544_wire_constant <= "11101000";
    type_cast_5546_wire_constant <= "00110111";
    type_cast_5554_wire_constant <= "01110101";
    type_cast_5556_wire_constant <= "00011100";
    type_cast_5564_wire_constant <= "01101110";
    type_cast_5566_wire_constant <= "11011111";
    type_cast_5574_wire_constant <= "11110001";
    type_cast_5576_wire_constant <= "01000111";
    type_cast_5584_wire_constant <= "01110001";
    type_cast_5586_wire_constant <= "00011010";
    type_cast_5594_wire_constant <= "00101001";
    type_cast_5596_wire_constant <= "00011101";
    type_cast_5604_wire_constant <= "10001001";
    type_cast_5606_wire_constant <= "11000101";
    type_cast_5614_wire_constant <= "10110111";
    type_cast_5616_wire_constant <= "01101111";
    type_cast_5624_wire_constant <= "00001110";
    type_cast_5626_wire_constant <= "01100010";
    type_cast_5634_wire_constant <= "00011000";
    type_cast_5636_wire_constant <= "10101010";
    type_cast_5644_wire_constant <= "00011011";
    type_cast_5646_wire_constant <= "10111110";
    type_cast_5654_wire_constant <= "01010110";
    type_cast_5656_wire_constant <= "11111100";
    type_cast_5664_wire_constant <= "01001011";
    type_cast_5666_wire_constant <= "00111110";
    type_cast_5674_wire_constant <= "11010010";
    type_cast_5676_wire_constant <= "11000110";
    type_cast_5684_wire_constant <= "00100000";
    type_cast_5686_wire_constant <= "01111001";
    type_cast_5694_wire_constant <= "11011011";
    type_cast_5696_wire_constant <= "10011010";
    type_cast_5704_wire_constant <= "11111110";
    type_cast_5706_wire_constant <= "11000000";
    type_cast_5714_wire_constant <= "11001101";
    type_cast_5716_wire_constant <= "01111000";
    type_cast_5724_wire_constant <= "11110100";
    type_cast_5726_wire_constant <= "01011010";
    type_cast_5734_wire_constant <= "11011101";
    type_cast_5736_wire_constant <= "00011111";
    type_cast_5744_wire_constant <= "00110011";
    type_cast_5746_wire_constant <= "10101000";
    type_cast_5754_wire_constant <= "00000111";
    type_cast_5756_wire_constant <= "10001000";
    type_cast_5764_wire_constant <= "00110001";
    type_cast_5766_wire_constant <= "11000111";
    type_cast_5774_wire_constant <= "00010010";
    type_cast_5776_wire_constant <= "10110001";
    type_cast_5784_wire_constant <= "01011001";
    type_cast_5786_wire_constant <= "00010000";
    type_cast_5794_wire_constant <= "10000000";
    type_cast_5796_wire_constant <= "00100111";
    type_cast_5804_wire_constant <= "01011111";
    type_cast_5806_wire_constant <= "11101100";
    type_cast_5814_wire_constant <= "01010001";
    type_cast_5816_wire_constant <= "01100000";
    type_cast_5824_wire_constant <= "10101001";
    type_cast_5826_wire_constant <= "01111111";
    type_cast_5834_wire_constant <= "10110101";
    type_cast_5836_wire_constant <= "00011001";
    type_cast_5844_wire_constant <= "00001101";
    type_cast_5846_wire_constant <= "01001010";
    type_cast_5854_wire_constant <= "11100101";
    type_cast_5856_wire_constant <= "00101101";
    type_cast_5864_wire_constant <= "10011111";
    type_cast_5866_wire_constant <= "01111010";
    type_cast_5874_wire_constant <= "11001001";
    type_cast_5876_wire_constant <= "10010011";
    type_cast_5884_wire_constant <= "11101111";
    type_cast_5886_wire_constant <= "10011100";
    type_cast_5894_wire_constant <= "11100000";
    type_cast_5896_wire_constant <= "10100000";
    type_cast_5904_wire_constant <= "01001101";
    type_cast_5906_wire_constant <= "00111011";
    type_cast_5914_wire_constant <= "00101010";
    type_cast_5916_wire_constant <= "10101110";
    type_cast_5924_wire_constant <= "10110000";
    type_cast_5926_wire_constant <= "11110101";
    type_cast_5934_wire_constant <= "11101011";
    type_cast_5936_wire_constant <= "11001000";
    type_cast_5944_wire_constant <= "00111100";
    type_cast_5946_wire_constant <= "10111011";
    type_cast_5954_wire_constant <= "01010011";
    type_cast_5956_wire_constant <= "10000011";
    type_cast_5964_wire_constant <= "01100001";
    type_cast_5966_wire_constant <= "10011001";
    type_cast_5974_wire_constant <= "00101011";
    type_cast_5976_wire_constant <= "00010111";
    type_cast_5984_wire_constant <= "01111110";
    type_cast_5986_wire_constant <= "00000100";
    type_cast_5994_wire_constant <= "01110111";
    type_cast_5996_wire_constant <= "10111010";
    type_cast_6004_wire_constant <= "00100110";
    type_cast_6006_wire_constant <= "11010110";
    type_cast_6014_wire_constant <= "01101001";
    type_cast_6016_wire_constant <= "11100001";
    type_cast_6024_wire_constant <= "01100011";
    type_cast_6026_wire_constant <= "00010100";
    type_cast_6034_wire_constant <= "00100001";
    type_cast_6036_wire_constant <= "01010101";
    type_cast_6044_wire_constant <= "01111101";
    type_cast_6046_wire_constant <= "00001100";
    -- flow-through select operator MUX_4777_inst
    IMA0_4778 <= type_cast_4774_wire_constant when (BITSEL_u8_u1_4772_wire(0) /=  '0') else type_cast_4776_wire_constant;
    -- flow-through select operator MUX_4787_inst
    IMA1_4788 <= type_cast_4784_wire_constant when (BITSEL_u8_u1_4782_wire(0) /=  '0') else type_cast_4786_wire_constant;
    -- flow-through select operator MUX_4797_inst
    IMA2_4798 <= type_cast_4794_wire_constant when (BITSEL_u8_u1_4792_wire(0) /=  '0') else type_cast_4796_wire_constant;
    -- flow-through select operator MUX_4807_inst
    IMA3_4808 <= type_cast_4804_wire_constant when (BITSEL_u8_u1_4802_wire(0) /=  '0') else type_cast_4806_wire_constant;
    -- flow-through select operator MUX_4817_inst
    IMA4_4818 <= type_cast_4814_wire_constant when (BITSEL_u8_u1_4812_wire(0) /=  '0') else type_cast_4816_wire_constant;
    -- flow-through select operator MUX_4827_inst
    IMA5_4828 <= type_cast_4824_wire_constant when (BITSEL_u8_u1_4822_wire(0) /=  '0') else type_cast_4826_wire_constant;
    -- flow-through select operator MUX_4837_inst
    IMA6_4838 <= type_cast_4834_wire_constant when (BITSEL_u8_u1_4832_wire(0) /=  '0') else type_cast_4836_wire_constant;
    -- flow-through select operator MUX_4847_inst
    IMA7_4848 <= type_cast_4844_wire_constant when (BITSEL_u8_u1_4842_wire(0) /=  '0') else type_cast_4846_wire_constant;
    -- flow-through select operator MUX_4857_inst
    IMA8_4858 <= type_cast_4854_wire_constant when (BITSEL_u8_u1_4852_wire(0) /=  '0') else type_cast_4856_wire_constant;
    -- flow-through select operator MUX_4867_inst
    IMA9_4868 <= type_cast_4864_wire_constant when (BITSEL_u8_u1_4862_wire(0) /=  '0') else type_cast_4866_wire_constant;
    -- flow-through select operator MUX_4877_inst
    IMA10_4878 <= type_cast_4874_wire_constant when (BITSEL_u8_u1_4872_wire(0) /=  '0') else type_cast_4876_wire_constant;
    -- flow-through select operator MUX_4887_inst
    IMA11_4888 <= type_cast_4884_wire_constant when (BITSEL_u8_u1_4882_wire(0) /=  '0') else type_cast_4886_wire_constant;
    -- flow-through select operator MUX_4897_inst
    IMA12_4898 <= type_cast_4894_wire_constant when (BITSEL_u8_u1_4892_wire(0) /=  '0') else type_cast_4896_wire_constant;
    -- flow-through select operator MUX_4907_inst
    IMA13_4908 <= type_cast_4904_wire_constant when (BITSEL_u8_u1_4902_wire(0) /=  '0') else type_cast_4906_wire_constant;
    -- flow-through select operator MUX_4917_inst
    IMA14_4918 <= type_cast_4914_wire_constant when (BITSEL_u8_u1_4912_wire(0) /=  '0') else type_cast_4916_wire_constant;
    -- flow-through select operator MUX_4927_inst
    IMA15_4928 <= type_cast_4924_wire_constant when (BITSEL_u8_u1_4922_wire(0) /=  '0') else type_cast_4926_wire_constant;
    -- flow-through select operator MUX_4937_inst
    IMA16_4938 <= type_cast_4934_wire_constant when (BITSEL_u8_u1_4932_wire(0) /=  '0') else type_cast_4936_wire_constant;
    -- flow-through select operator MUX_4947_inst
    IMA17_4948 <= type_cast_4944_wire_constant when (BITSEL_u8_u1_4942_wire(0) /=  '0') else type_cast_4946_wire_constant;
    -- flow-through select operator MUX_4957_inst
    IMA18_4958 <= type_cast_4954_wire_constant when (BITSEL_u8_u1_4952_wire(0) /=  '0') else type_cast_4956_wire_constant;
    -- flow-through select operator MUX_4967_inst
    IMA19_4968 <= type_cast_4964_wire_constant when (BITSEL_u8_u1_4962_wire(0) /=  '0') else type_cast_4966_wire_constant;
    -- flow-through select operator MUX_4977_inst
    IMA20_4978 <= type_cast_4974_wire_constant when (BITSEL_u8_u1_4972_wire(0) /=  '0') else type_cast_4976_wire_constant;
    -- flow-through select operator MUX_4987_inst
    IMA21_4988 <= type_cast_4984_wire_constant when (BITSEL_u8_u1_4982_wire(0) /=  '0') else type_cast_4986_wire_constant;
    -- flow-through select operator MUX_4997_inst
    IMA22_4998 <= type_cast_4994_wire_constant when (BITSEL_u8_u1_4992_wire(0) /=  '0') else type_cast_4996_wire_constant;
    -- flow-through select operator MUX_5007_inst
    IMA23_5008 <= type_cast_5004_wire_constant when (BITSEL_u8_u1_5002_wire(0) /=  '0') else type_cast_5006_wire_constant;
    -- flow-through select operator MUX_5017_inst
    IMA24_5018 <= type_cast_5014_wire_constant when (BITSEL_u8_u1_5012_wire(0) /=  '0') else type_cast_5016_wire_constant;
    -- flow-through select operator MUX_5027_inst
    IMA25_5028 <= type_cast_5024_wire_constant when (BITSEL_u8_u1_5022_wire(0) /=  '0') else type_cast_5026_wire_constant;
    -- flow-through select operator MUX_5037_inst
    IMA26_5038 <= type_cast_5034_wire_constant when (BITSEL_u8_u1_5032_wire(0) /=  '0') else type_cast_5036_wire_constant;
    -- flow-through select operator MUX_5047_inst
    IMA27_5048 <= type_cast_5044_wire_constant when (BITSEL_u8_u1_5042_wire(0) /=  '0') else type_cast_5046_wire_constant;
    -- flow-through select operator MUX_5057_inst
    IMA28_5058 <= type_cast_5054_wire_constant when (BITSEL_u8_u1_5052_wire(0) /=  '0') else type_cast_5056_wire_constant;
    -- flow-through select operator MUX_5067_inst
    IMA29_5068 <= type_cast_5064_wire_constant when (BITSEL_u8_u1_5062_wire(0) /=  '0') else type_cast_5066_wire_constant;
    -- flow-through select operator MUX_5077_inst
    IMA30_5078 <= type_cast_5074_wire_constant when (BITSEL_u8_u1_5072_wire(0) /=  '0') else type_cast_5076_wire_constant;
    -- flow-through select operator MUX_5087_inst
    IMA31_5088 <= type_cast_5084_wire_constant when (BITSEL_u8_u1_5082_wire(0) /=  '0') else type_cast_5086_wire_constant;
    -- flow-through select operator MUX_5097_inst
    IMA32_5098 <= type_cast_5094_wire_constant when (BITSEL_u8_u1_5092_wire(0) /=  '0') else type_cast_5096_wire_constant;
    -- flow-through select operator MUX_5107_inst
    IMA33_5108 <= type_cast_5104_wire_constant when (BITSEL_u8_u1_5102_wire(0) /=  '0') else type_cast_5106_wire_constant;
    -- flow-through select operator MUX_5117_inst
    IMA34_5118 <= type_cast_5114_wire_constant when (BITSEL_u8_u1_5112_wire(0) /=  '0') else type_cast_5116_wire_constant;
    -- flow-through select operator MUX_5127_inst
    IMA35_5128 <= type_cast_5124_wire_constant when (BITSEL_u8_u1_5122_wire(0) /=  '0') else type_cast_5126_wire_constant;
    -- flow-through select operator MUX_5137_inst
    IMA36_5138 <= type_cast_5134_wire_constant when (BITSEL_u8_u1_5132_wire(0) /=  '0') else type_cast_5136_wire_constant;
    -- flow-through select operator MUX_5147_inst
    IMA37_5148 <= type_cast_5144_wire_constant when (BITSEL_u8_u1_5142_wire(0) /=  '0') else type_cast_5146_wire_constant;
    -- flow-through select operator MUX_5157_inst
    IMA38_5158 <= type_cast_5154_wire_constant when (BITSEL_u8_u1_5152_wire(0) /=  '0') else type_cast_5156_wire_constant;
    -- flow-through select operator MUX_5167_inst
    IMA39_5168 <= type_cast_5164_wire_constant when (BITSEL_u8_u1_5162_wire(0) /=  '0') else type_cast_5166_wire_constant;
    -- flow-through select operator MUX_5177_inst
    IMA40_5178 <= type_cast_5174_wire_constant when (BITSEL_u8_u1_5172_wire(0) /=  '0') else type_cast_5176_wire_constant;
    -- flow-through select operator MUX_5187_inst
    IMA41_5188 <= type_cast_5184_wire_constant when (BITSEL_u8_u1_5182_wire(0) /=  '0') else type_cast_5186_wire_constant;
    -- flow-through select operator MUX_5197_inst
    IMA42_5198 <= type_cast_5194_wire_constant when (BITSEL_u8_u1_5192_wire(0) /=  '0') else type_cast_5196_wire_constant;
    -- flow-through select operator MUX_5207_inst
    IMA43_5208 <= type_cast_5204_wire_constant when (BITSEL_u8_u1_5202_wire(0) /=  '0') else type_cast_5206_wire_constant;
    -- flow-through select operator MUX_5217_inst
    IMA44_5218 <= type_cast_5214_wire_constant when (BITSEL_u8_u1_5212_wire(0) /=  '0') else type_cast_5216_wire_constant;
    -- flow-through select operator MUX_5227_inst
    IMA45_5228 <= type_cast_5224_wire_constant when (BITSEL_u8_u1_5222_wire(0) /=  '0') else type_cast_5226_wire_constant;
    -- flow-through select operator MUX_5237_inst
    IMA46_5238 <= type_cast_5234_wire_constant when (BITSEL_u8_u1_5232_wire(0) /=  '0') else type_cast_5236_wire_constant;
    -- flow-through select operator MUX_5247_inst
    IMA47_5248 <= type_cast_5244_wire_constant when (BITSEL_u8_u1_5242_wire(0) /=  '0') else type_cast_5246_wire_constant;
    -- flow-through select operator MUX_5257_inst
    IMA48_5258 <= type_cast_5254_wire_constant when (BITSEL_u8_u1_5252_wire(0) /=  '0') else type_cast_5256_wire_constant;
    -- flow-through select operator MUX_5267_inst
    IMA49_5268 <= type_cast_5264_wire_constant when (BITSEL_u8_u1_5262_wire(0) /=  '0') else type_cast_5266_wire_constant;
    -- flow-through select operator MUX_5277_inst
    IMA50_5278 <= type_cast_5274_wire_constant when (BITSEL_u8_u1_5272_wire(0) /=  '0') else type_cast_5276_wire_constant;
    -- flow-through select operator MUX_5287_inst
    IMA51_5288 <= type_cast_5284_wire_constant when (BITSEL_u8_u1_5282_wire(0) /=  '0') else type_cast_5286_wire_constant;
    -- flow-through select operator MUX_5297_inst
    IMA52_5298 <= type_cast_5294_wire_constant when (BITSEL_u8_u1_5292_wire(0) /=  '0') else type_cast_5296_wire_constant;
    -- flow-through select operator MUX_5307_inst
    IMA53_5308 <= type_cast_5304_wire_constant when (BITSEL_u8_u1_5302_wire(0) /=  '0') else type_cast_5306_wire_constant;
    -- flow-through select operator MUX_5317_inst
    IMA54_5318 <= type_cast_5314_wire_constant when (BITSEL_u8_u1_5312_wire(0) /=  '0') else type_cast_5316_wire_constant;
    -- flow-through select operator MUX_5327_inst
    IMA55_5328 <= type_cast_5324_wire_constant when (BITSEL_u8_u1_5322_wire(0) /=  '0') else type_cast_5326_wire_constant;
    -- flow-through select operator MUX_5337_inst
    IMA56_5338 <= type_cast_5334_wire_constant when (BITSEL_u8_u1_5332_wire(0) /=  '0') else type_cast_5336_wire_constant;
    -- flow-through select operator MUX_5347_inst
    IMA57_5348 <= type_cast_5344_wire_constant when (BITSEL_u8_u1_5342_wire(0) /=  '0') else type_cast_5346_wire_constant;
    -- flow-through select operator MUX_5357_inst
    IMA58_5358 <= type_cast_5354_wire_constant when (BITSEL_u8_u1_5352_wire(0) /=  '0') else type_cast_5356_wire_constant;
    -- flow-through select operator MUX_5367_inst
    IMA59_5368 <= type_cast_5364_wire_constant when (BITSEL_u8_u1_5362_wire(0) /=  '0') else type_cast_5366_wire_constant;
    -- flow-through select operator MUX_5377_inst
    IMA60_5378 <= type_cast_5374_wire_constant when (BITSEL_u8_u1_5372_wire(0) /=  '0') else type_cast_5376_wire_constant;
    -- flow-through select operator MUX_5387_inst
    IMA61_5388 <= type_cast_5384_wire_constant when (BITSEL_u8_u1_5382_wire(0) /=  '0') else type_cast_5386_wire_constant;
    -- flow-through select operator MUX_5397_inst
    IMA62_5398 <= type_cast_5394_wire_constant when (BITSEL_u8_u1_5392_wire(0) /=  '0') else type_cast_5396_wire_constant;
    -- flow-through select operator MUX_5407_inst
    IMA63_5408 <= type_cast_5404_wire_constant when (BITSEL_u8_u1_5402_wire(0) /=  '0') else type_cast_5406_wire_constant;
    -- flow-through select operator MUX_5417_inst
    IMA64_5418 <= type_cast_5414_wire_constant when (BITSEL_u8_u1_5412_wire(0) /=  '0') else type_cast_5416_wire_constant;
    -- flow-through select operator MUX_5427_inst
    IMA65_5428 <= type_cast_5424_wire_constant when (BITSEL_u8_u1_5422_wire(0) /=  '0') else type_cast_5426_wire_constant;
    -- flow-through select operator MUX_5437_inst
    IMA66_5438 <= type_cast_5434_wire_constant when (BITSEL_u8_u1_5432_wire(0) /=  '0') else type_cast_5436_wire_constant;
    -- flow-through select operator MUX_5447_inst
    IMA67_5448 <= type_cast_5444_wire_constant when (BITSEL_u8_u1_5442_wire(0) /=  '0') else type_cast_5446_wire_constant;
    -- flow-through select operator MUX_5457_inst
    IMA68_5458 <= type_cast_5454_wire_constant when (BITSEL_u8_u1_5452_wire(0) /=  '0') else type_cast_5456_wire_constant;
    -- flow-through select operator MUX_5467_inst
    IMA69_5468 <= type_cast_5464_wire_constant when (BITSEL_u8_u1_5462_wire(0) /=  '0') else type_cast_5466_wire_constant;
    -- flow-through select operator MUX_5477_inst
    IMA70_5478 <= type_cast_5474_wire_constant when (BITSEL_u8_u1_5472_wire(0) /=  '0') else type_cast_5476_wire_constant;
    -- flow-through select operator MUX_5487_inst
    IMA71_5488 <= type_cast_5484_wire_constant when (BITSEL_u8_u1_5482_wire(0) /=  '0') else type_cast_5486_wire_constant;
    -- flow-through select operator MUX_5497_inst
    IMA72_5498 <= type_cast_5494_wire_constant when (BITSEL_u8_u1_5492_wire(0) /=  '0') else type_cast_5496_wire_constant;
    -- flow-through select operator MUX_5507_inst
    IMA73_5508 <= type_cast_5504_wire_constant when (BITSEL_u8_u1_5502_wire(0) /=  '0') else type_cast_5506_wire_constant;
    -- flow-through select operator MUX_5517_inst
    IMA74_5518 <= type_cast_5514_wire_constant when (BITSEL_u8_u1_5512_wire(0) /=  '0') else type_cast_5516_wire_constant;
    -- flow-through select operator MUX_5527_inst
    IMA75_5528 <= type_cast_5524_wire_constant when (BITSEL_u8_u1_5522_wire(0) /=  '0') else type_cast_5526_wire_constant;
    -- flow-through select operator MUX_5537_inst
    IMA76_5538 <= type_cast_5534_wire_constant when (BITSEL_u8_u1_5532_wire(0) /=  '0') else type_cast_5536_wire_constant;
    -- flow-through select operator MUX_5547_inst
    IMA77_5548 <= type_cast_5544_wire_constant when (BITSEL_u8_u1_5542_wire(0) /=  '0') else type_cast_5546_wire_constant;
    -- flow-through select operator MUX_5557_inst
    IMA78_5558 <= type_cast_5554_wire_constant when (BITSEL_u8_u1_5552_wire(0) /=  '0') else type_cast_5556_wire_constant;
    -- flow-through select operator MUX_5567_inst
    IMA79_5568 <= type_cast_5564_wire_constant when (BITSEL_u8_u1_5562_wire(0) /=  '0') else type_cast_5566_wire_constant;
    -- flow-through select operator MUX_5577_inst
    IMA80_5578 <= type_cast_5574_wire_constant when (BITSEL_u8_u1_5572_wire(0) /=  '0') else type_cast_5576_wire_constant;
    -- flow-through select operator MUX_5587_inst
    IMA81_5588 <= type_cast_5584_wire_constant when (BITSEL_u8_u1_5582_wire(0) /=  '0') else type_cast_5586_wire_constant;
    -- flow-through select operator MUX_5597_inst
    IMA82_5598 <= type_cast_5594_wire_constant when (BITSEL_u8_u1_5592_wire(0) /=  '0') else type_cast_5596_wire_constant;
    -- flow-through select operator MUX_5607_inst
    IMA83_5608 <= type_cast_5604_wire_constant when (BITSEL_u8_u1_5602_wire(0) /=  '0') else type_cast_5606_wire_constant;
    -- flow-through select operator MUX_5617_inst
    IMA84_5618 <= type_cast_5614_wire_constant when (BITSEL_u8_u1_5612_wire(0) /=  '0') else type_cast_5616_wire_constant;
    -- flow-through select operator MUX_5627_inst
    IMA85_5628 <= type_cast_5624_wire_constant when (BITSEL_u8_u1_5622_wire(0) /=  '0') else type_cast_5626_wire_constant;
    -- flow-through select operator MUX_5637_inst
    IMA86_5638 <= type_cast_5634_wire_constant when (BITSEL_u8_u1_5632_wire(0) /=  '0') else type_cast_5636_wire_constant;
    -- flow-through select operator MUX_5647_inst
    IMA87_5648 <= type_cast_5644_wire_constant when (BITSEL_u8_u1_5642_wire(0) /=  '0') else type_cast_5646_wire_constant;
    -- flow-through select operator MUX_5657_inst
    IMA88_5658 <= type_cast_5654_wire_constant when (BITSEL_u8_u1_5652_wire(0) /=  '0') else type_cast_5656_wire_constant;
    -- flow-through select operator MUX_5667_inst
    IMA89_5668 <= type_cast_5664_wire_constant when (BITSEL_u8_u1_5662_wire(0) /=  '0') else type_cast_5666_wire_constant;
    -- flow-through select operator MUX_5677_inst
    IMA90_5678 <= type_cast_5674_wire_constant when (BITSEL_u8_u1_5672_wire(0) /=  '0') else type_cast_5676_wire_constant;
    -- flow-through select operator MUX_5687_inst
    IMA91_5688 <= type_cast_5684_wire_constant when (BITSEL_u8_u1_5682_wire(0) /=  '0') else type_cast_5686_wire_constant;
    -- flow-through select operator MUX_5697_inst
    IMA92_5698 <= type_cast_5694_wire_constant when (BITSEL_u8_u1_5692_wire(0) /=  '0') else type_cast_5696_wire_constant;
    -- flow-through select operator MUX_5707_inst
    IMA93_5708 <= type_cast_5704_wire_constant when (BITSEL_u8_u1_5702_wire(0) /=  '0') else type_cast_5706_wire_constant;
    -- flow-through select operator MUX_5717_inst
    IMA94_5718 <= type_cast_5714_wire_constant when (BITSEL_u8_u1_5712_wire(0) /=  '0') else type_cast_5716_wire_constant;
    -- flow-through select operator MUX_5727_inst
    IMA95_5728 <= type_cast_5724_wire_constant when (BITSEL_u8_u1_5722_wire(0) /=  '0') else type_cast_5726_wire_constant;
    -- flow-through select operator MUX_5737_inst
    IMA96_5738 <= type_cast_5734_wire_constant when (BITSEL_u8_u1_5732_wire(0) /=  '0') else type_cast_5736_wire_constant;
    -- flow-through select operator MUX_5747_inst
    IMA97_5748 <= type_cast_5744_wire_constant when (BITSEL_u8_u1_5742_wire(0) /=  '0') else type_cast_5746_wire_constant;
    -- flow-through select operator MUX_5757_inst
    IMA98_5758 <= type_cast_5754_wire_constant when (BITSEL_u8_u1_5752_wire(0) /=  '0') else type_cast_5756_wire_constant;
    -- flow-through select operator MUX_5767_inst
    IMA99_5768 <= type_cast_5764_wire_constant when (BITSEL_u8_u1_5762_wire(0) /=  '0') else type_cast_5766_wire_constant;
    -- flow-through select operator MUX_5777_inst
    IMA100_5778 <= type_cast_5774_wire_constant when (BITSEL_u8_u1_5772_wire(0) /=  '0') else type_cast_5776_wire_constant;
    -- flow-through select operator MUX_5787_inst
    IMA101_5788 <= type_cast_5784_wire_constant when (BITSEL_u8_u1_5782_wire(0) /=  '0') else type_cast_5786_wire_constant;
    -- flow-through select operator MUX_5797_inst
    IMA102_5798 <= type_cast_5794_wire_constant when (BITSEL_u8_u1_5792_wire(0) /=  '0') else type_cast_5796_wire_constant;
    -- flow-through select operator MUX_5807_inst
    IMA103_5808 <= type_cast_5804_wire_constant when (BITSEL_u8_u1_5802_wire(0) /=  '0') else type_cast_5806_wire_constant;
    -- flow-through select operator MUX_5817_inst
    IMA104_5818 <= type_cast_5814_wire_constant when (BITSEL_u8_u1_5812_wire(0) /=  '0') else type_cast_5816_wire_constant;
    -- flow-through select operator MUX_5827_inst
    IMA105_5828 <= type_cast_5824_wire_constant when (BITSEL_u8_u1_5822_wire(0) /=  '0') else type_cast_5826_wire_constant;
    -- flow-through select operator MUX_5837_inst
    IMA106_5838 <= type_cast_5834_wire_constant when (BITSEL_u8_u1_5832_wire(0) /=  '0') else type_cast_5836_wire_constant;
    -- flow-through select operator MUX_5847_inst
    IMA107_5848 <= type_cast_5844_wire_constant when (BITSEL_u8_u1_5842_wire(0) /=  '0') else type_cast_5846_wire_constant;
    -- flow-through select operator MUX_5857_inst
    IMA108_5858 <= type_cast_5854_wire_constant when (BITSEL_u8_u1_5852_wire(0) /=  '0') else type_cast_5856_wire_constant;
    -- flow-through select operator MUX_5867_inst
    IMA109_5868 <= type_cast_5864_wire_constant when (BITSEL_u8_u1_5862_wire(0) /=  '0') else type_cast_5866_wire_constant;
    -- flow-through select operator MUX_5877_inst
    IMA110_5878 <= type_cast_5874_wire_constant when (BITSEL_u8_u1_5872_wire(0) /=  '0') else type_cast_5876_wire_constant;
    -- flow-through select operator MUX_5887_inst
    IMA111_5888 <= type_cast_5884_wire_constant when (BITSEL_u8_u1_5882_wire(0) /=  '0') else type_cast_5886_wire_constant;
    -- flow-through select operator MUX_5897_inst
    IMA112_5898 <= type_cast_5894_wire_constant when (BITSEL_u8_u1_5892_wire(0) /=  '0') else type_cast_5896_wire_constant;
    -- flow-through select operator MUX_5907_inst
    IMA113_5908 <= type_cast_5904_wire_constant when (BITSEL_u8_u1_5902_wire(0) /=  '0') else type_cast_5906_wire_constant;
    -- flow-through select operator MUX_5917_inst
    IMA114_5918 <= type_cast_5914_wire_constant when (BITSEL_u8_u1_5912_wire(0) /=  '0') else type_cast_5916_wire_constant;
    -- flow-through select operator MUX_5927_inst
    IMA115_5928 <= type_cast_5924_wire_constant when (BITSEL_u8_u1_5922_wire(0) /=  '0') else type_cast_5926_wire_constant;
    -- flow-through select operator MUX_5937_inst
    IMA116_5938 <= type_cast_5934_wire_constant when (BITSEL_u8_u1_5932_wire(0) /=  '0') else type_cast_5936_wire_constant;
    -- flow-through select operator MUX_5947_inst
    IMA117_5948 <= type_cast_5944_wire_constant when (BITSEL_u8_u1_5942_wire(0) /=  '0') else type_cast_5946_wire_constant;
    -- flow-through select operator MUX_5957_inst
    IMA118_5958 <= type_cast_5954_wire_constant when (BITSEL_u8_u1_5952_wire(0) /=  '0') else type_cast_5956_wire_constant;
    -- flow-through select operator MUX_5967_inst
    IMA119_5968 <= type_cast_5964_wire_constant when (BITSEL_u8_u1_5962_wire(0) /=  '0') else type_cast_5966_wire_constant;
    -- flow-through select operator MUX_5977_inst
    IMA120_5978 <= type_cast_5974_wire_constant when (BITSEL_u8_u1_5972_wire(0) /=  '0') else type_cast_5976_wire_constant;
    -- flow-through select operator MUX_5987_inst
    IMA121_5988 <= type_cast_5984_wire_constant when (BITSEL_u8_u1_5982_wire(0) /=  '0') else type_cast_5986_wire_constant;
    -- flow-through select operator MUX_5997_inst
    IMA122_5998 <= type_cast_5994_wire_constant when (BITSEL_u8_u1_5992_wire(0) /=  '0') else type_cast_5996_wire_constant;
    -- flow-through select operator MUX_6007_inst
    IMA123_6008 <= type_cast_6004_wire_constant when (BITSEL_u8_u1_6002_wire(0) /=  '0') else type_cast_6006_wire_constant;
    -- flow-through select operator MUX_6017_inst
    IMA124_6018 <= type_cast_6014_wire_constant when (BITSEL_u8_u1_6012_wire(0) /=  '0') else type_cast_6016_wire_constant;
    -- flow-through select operator MUX_6027_inst
    IMA125_6028 <= type_cast_6024_wire_constant when (BITSEL_u8_u1_6022_wire(0) /=  '0') else type_cast_6026_wire_constant;
    -- flow-through select operator MUX_6037_inst
    IMA126_6038 <= type_cast_6034_wire_constant when (BITSEL_u8_u1_6032_wire(0) /=  '0') else type_cast_6036_wire_constant;
    -- flow-through select operator MUX_6047_inst
    IMA127_6048 <= type_cast_6044_wire_constant when (BITSEL_u8_u1_6042_wire(0) /=  '0') else type_cast_6046_wire_constant;
    -- flow-through select operator MUX_6055_inst
    IMB0_6056 <= IMA1_4788 when (BITSEL_u8_u1_6052_wire(0) /=  '0') else IMA0_4778;
    -- flow-through select operator MUX_6063_inst
    IMB1_6064 <= IMA3_4808 when (BITSEL_u8_u1_6060_wire(0) /=  '0') else IMA2_4798;
    -- flow-through select operator MUX_6071_inst
    IMB2_6072 <= IMA5_4828 when (BITSEL_u8_u1_6068_wire(0) /=  '0') else IMA4_4818;
    -- flow-through select operator MUX_6079_inst
    IMB3_6080 <= IMA7_4848 when (BITSEL_u8_u1_6076_wire(0) /=  '0') else IMA6_4838;
    -- flow-through select operator MUX_6087_inst
    IMB4_6088 <= IMA9_4868 when (BITSEL_u8_u1_6084_wire(0) /=  '0') else IMA8_4858;
    -- flow-through select operator MUX_6095_inst
    IMB5_6096 <= IMA11_4888 when (BITSEL_u8_u1_6092_wire(0) /=  '0') else IMA10_4878;
    -- flow-through select operator MUX_6103_inst
    IMB6_6104 <= IMA13_4908 when (BITSEL_u8_u1_6100_wire(0) /=  '0') else IMA12_4898;
    -- flow-through select operator MUX_6111_inst
    IMB7_6112 <= IMA15_4928 when (BITSEL_u8_u1_6108_wire(0) /=  '0') else IMA14_4918;
    -- flow-through select operator MUX_6119_inst
    IMB8_6120 <= IMA17_4948 when (BITSEL_u8_u1_6116_wire(0) /=  '0') else IMA16_4938;
    -- flow-through select operator MUX_6127_inst
    IMB9_6128 <= IMA19_4968 when (BITSEL_u8_u1_6124_wire(0) /=  '0') else IMA18_4958;
    -- flow-through select operator MUX_6135_inst
    IMB10_6136 <= IMA21_4988 when (BITSEL_u8_u1_6132_wire(0) /=  '0') else IMA20_4978;
    -- flow-through select operator MUX_6143_inst
    IMB11_6144 <= IMA23_5008 when (BITSEL_u8_u1_6140_wire(0) /=  '0') else IMA22_4998;
    -- flow-through select operator MUX_6151_inst
    IMB12_6152 <= IMA25_5028 when (BITSEL_u8_u1_6148_wire(0) /=  '0') else IMA24_5018;
    -- flow-through select operator MUX_6159_inst
    IMB13_6160 <= IMA27_5048 when (BITSEL_u8_u1_6156_wire(0) /=  '0') else IMA26_5038;
    -- flow-through select operator MUX_6167_inst
    IMB14_6168 <= IMA29_5068 when (BITSEL_u8_u1_6164_wire(0) /=  '0') else IMA28_5058;
    -- flow-through select operator MUX_6175_inst
    IMB15_6176 <= IMA31_5088 when (BITSEL_u8_u1_6172_wire(0) /=  '0') else IMA30_5078;
    -- flow-through select operator MUX_6183_inst
    IMB16_6184 <= IMA33_5108 when (BITSEL_u8_u1_6180_wire(0) /=  '0') else IMA32_5098;
    -- flow-through select operator MUX_6191_inst
    IMB17_6192 <= IMA35_5128 when (BITSEL_u8_u1_6188_wire(0) /=  '0') else IMA34_5118;
    -- flow-through select operator MUX_6199_inst
    IMB18_6200 <= IMA37_5148 when (BITSEL_u8_u1_6196_wire(0) /=  '0') else IMA36_5138;
    -- flow-through select operator MUX_6207_inst
    IMB19_6208 <= IMA39_5168 when (BITSEL_u8_u1_6204_wire(0) /=  '0') else IMA38_5158;
    -- flow-through select operator MUX_6215_inst
    IMB20_6216 <= IMA41_5188 when (BITSEL_u8_u1_6212_wire(0) /=  '0') else IMA40_5178;
    -- flow-through select operator MUX_6223_inst
    IMB21_6224 <= IMA43_5208 when (BITSEL_u8_u1_6220_wire(0) /=  '0') else IMA42_5198;
    -- flow-through select operator MUX_6231_inst
    IMB22_6232 <= IMA45_5228 when (BITSEL_u8_u1_6228_wire(0) /=  '0') else IMA44_5218;
    -- flow-through select operator MUX_6239_inst
    IMB23_6240 <= IMA47_5248 when (BITSEL_u8_u1_6236_wire(0) /=  '0') else IMA46_5238;
    -- flow-through select operator MUX_6247_inst
    IMB24_6248 <= IMA49_5268 when (BITSEL_u8_u1_6244_wire(0) /=  '0') else IMA48_5258;
    -- flow-through select operator MUX_6255_inst
    IMB25_6256 <= IMA51_5288 when (BITSEL_u8_u1_6252_wire(0) /=  '0') else IMA50_5278;
    -- flow-through select operator MUX_6263_inst
    IMB26_6264 <= IMA53_5308 when (BITSEL_u8_u1_6260_wire(0) /=  '0') else IMA52_5298;
    -- flow-through select operator MUX_6271_inst
    IMB27_6272 <= IMA55_5328 when (BITSEL_u8_u1_6268_wire(0) /=  '0') else IMA54_5318;
    -- flow-through select operator MUX_6279_inst
    IMB28_6280 <= IMA57_5348 when (BITSEL_u8_u1_6276_wire(0) /=  '0') else IMA56_5338;
    -- flow-through select operator MUX_6287_inst
    IMB29_6288 <= IMA59_5368 when (BITSEL_u8_u1_6284_wire(0) /=  '0') else IMA58_5358;
    -- flow-through select operator MUX_6295_inst
    IMB30_6296 <= IMA61_5388 when (BITSEL_u8_u1_6292_wire(0) /=  '0') else IMA60_5378;
    -- flow-through select operator MUX_6303_inst
    IMB31_6304 <= IMA63_5408 when (BITSEL_u8_u1_6300_wire(0) /=  '0') else IMA62_5398;
    -- flow-through select operator MUX_6311_inst
    IMB32_6312 <= IMA65_5428 when (BITSEL_u8_u1_6308_wire(0) /=  '0') else IMA64_5418;
    -- flow-through select operator MUX_6319_inst
    IMB33_6320 <= IMA67_5448 when (BITSEL_u8_u1_6316_wire(0) /=  '0') else IMA66_5438;
    -- flow-through select operator MUX_6327_inst
    IMB34_6328 <= IMA69_5468 when (BITSEL_u8_u1_6324_wire(0) /=  '0') else IMA68_5458;
    -- flow-through select operator MUX_6335_inst
    IMB35_6336 <= IMA71_5488 when (BITSEL_u8_u1_6332_wire(0) /=  '0') else IMA70_5478;
    -- flow-through select operator MUX_6343_inst
    IMB36_6344 <= IMA73_5508 when (BITSEL_u8_u1_6340_wire(0) /=  '0') else IMA72_5498;
    -- flow-through select operator MUX_6351_inst
    IMB37_6352 <= IMA75_5528 when (BITSEL_u8_u1_6348_wire(0) /=  '0') else IMA74_5518;
    -- flow-through select operator MUX_6359_inst
    IMB38_6360 <= IMA77_5548 when (BITSEL_u8_u1_6356_wire(0) /=  '0') else IMA76_5538;
    -- flow-through select operator MUX_6367_inst
    IMB39_6368 <= IMA79_5568 when (BITSEL_u8_u1_6364_wire(0) /=  '0') else IMA78_5558;
    -- flow-through select operator MUX_6375_inst
    IMB40_6376 <= IMA81_5588 when (BITSEL_u8_u1_6372_wire(0) /=  '0') else IMA80_5578;
    -- flow-through select operator MUX_6383_inst
    IMB41_6384 <= IMA83_5608 when (BITSEL_u8_u1_6380_wire(0) /=  '0') else IMA82_5598;
    -- flow-through select operator MUX_6391_inst
    IMB42_6392 <= IMA85_5628 when (BITSEL_u8_u1_6388_wire(0) /=  '0') else IMA84_5618;
    -- flow-through select operator MUX_6399_inst
    IMB43_6400 <= IMA87_5648 when (BITSEL_u8_u1_6396_wire(0) /=  '0') else IMA86_5638;
    -- flow-through select operator MUX_6407_inst
    IMB44_6408 <= IMA89_5668 when (BITSEL_u8_u1_6404_wire(0) /=  '0') else IMA88_5658;
    -- flow-through select operator MUX_6415_inst
    IMB45_6416 <= IMA91_5688 when (BITSEL_u8_u1_6412_wire(0) /=  '0') else IMA90_5678;
    -- flow-through select operator MUX_6423_inst
    IMB46_6424 <= IMA93_5708 when (BITSEL_u8_u1_6420_wire(0) /=  '0') else IMA92_5698;
    -- flow-through select operator MUX_6431_inst
    IMB47_6432 <= IMA95_5728 when (BITSEL_u8_u1_6428_wire(0) /=  '0') else IMA94_5718;
    -- flow-through select operator MUX_6439_inst
    IMB48_6440 <= IMA97_5748 when (BITSEL_u8_u1_6436_wire(0) /=  '0') else IMA96_5738;
    -- flow-through select operator MUX_6447_inst
    IMB49_6448 <= IMA99_5768 when (BITSEL_u8_u1_6444_wire(0) /=  '0') else IMA98_5758;
    -- flow-through select operator MUX_6455_inst
    IMB50_6456 <= IMA101_5788 when (BITSEL_u8_u1_6452_wire(0) /=  '0') else IMA100_5778;
    -- flow-through select operator MUX_6463_inst
    IMB51_6464 <= IMA103_5808 when (BITSEL_u8_u1_6460_wire(0) /=  '0') else IMA102_5798;
    -- flow-through select operator MUX_6471_inst
    IMB52_6472 <= IMA105_5828 when (BITSEL_u8_u1_6468_wire(0) /=  '0') else IMA104_5818;
    -- flow-through select operator MUX_6479_inst
    IMB53_6480 <= IMA107_5848 when (BITSEL_u8_u1_6476_wire(0) /=  '0') else IMA106_5838;
    -- flow-through select operator MUX_6487_inst
    IMB54_6488 <= IMA109_5868 when (BITSEL_u8_u1_6484_wire(0) /=  '0') else IMA108_5858;
    -- flow-through select operator MUX_6495_inst
    IMB55_6496 <= IMA111_5888 when (BITSEL_u8_u1_6492_wire(0) /=  '0') else IMA110_5878;
    -- flow-through select operator MUX_6503_inst
    IMB56_6504 <= IMA113_5908 when (BITSEL_u8_u1_6500_wire(0) /=  '0') else IMA112_5898;
    -- flow-through select operator MUX_6511_inst
    IMB57_6512 <= IMA115_5928 when (BITSEL_u8_u1_6508_wire(0) /=  '0') else IMA114_5918;
    -- flow-through select operator MUX_6519_inst
    IMB58_6520 <= IMA117_5948 when (BITSEL_u8_u1_6516_wire(0) /=  '0') else IMA116_5938;
    -- flow-through select operator MUX_6527_inst
    IMB59_6528 <= IMA119_5968 when (BITSEL_u8_u1_6524_wire(0) /=  '0') else IMA118_5958;
    -- flow-through select operator MUX_6535_inst
    IMB60_6536 <= IMA121_5988 when (BITSEL_u8_u1_6532_wire(0) /=  '0') else IMA120_5978;
    -- flow-through select operator MUX_6543_inst
    IMB61_6544 <= IMA123_6008 when (BITSEL_u8_u1_6540_wire(0) /=  '0') else IMA122_5998;
    -- flow-through select operator MUX_6551_inst
    IMB62_6552 <= IMA125_6028 when (BITSEL_u8_u1_6548_wire(0) /=  '0') else IMA124_6018;
    -- flow-through select operator MUX_6559_inst
    IMB63_6560 <= IMA127_6048 when (BITSEL_u8_u1_6556_wire(0) /=  '0') else IMA126_6038;
    -- flow-through select operator MUX_6567_inst
    IMC0_6568 <= IMB1_6064 when (BITSEL_u8_u1_6564_wire(0) /=  '0') else IMB0_6056;
    -- flow-through select operator MUX_6575_inst
    IMC1_6576 <= IMB3_6080 when (BITSEL_u8_u1_6572_wire(0) /=  '0') else IMB2_6072;
    -- flow-through select operator MUX_6583_inst
    IMC2_6584 <= IMB5_6096 when (BITSEL_u8_u1_6580_wire(0) /=  '0') else IMB4_6088;
    -- flow-through select operator MUX_6591_inst
    IMC3_6592 <= IMB7_6112 when (BITSEL_u8_u1_6588_wire(0) /=  '0') else IMB6_6104;
    -- flow-through select operator MUX_6599_inst
    IMC4_6600 <= IMB9_6128 when (BITSEL_u8_u1_6596_wire(0) /=  '0') else IMB8_6120;
    -- flow-through select operator MUX_6607_inst
    IMC5_6608 <= IMB11_6144 when (BITSEL_u8_u1_6604_wire(0) /=  '0') else IMB10_6136;
    -- flow-through select operator MUX_6615_inst
    IMC6_6616 <= IMB13_6160 when (BITSEL_u8_u1_6612_wire(0) /=  '0') else IMB12_6152;
    -- flow-through select operator MUX_6623_inst
    IMC7_6624 <= IMB15_6176 when (BITSEL_u8_u1_6620_wire(0) /=  '0') else IMB14_6168;
    -- flow-through select operator MUX_6631_inst
    IMC8_6632 <= IMB17_6192 when (BITSEL_u8_u1_6628_wire(0) /=  '0') else IMB16_6184;
    -- flow-through select operator MUX_6639_inst
    IMC9_6640 <= IMB19_6208 when (BITSEL_u8_u1_6636_wire(0) /=  '0') else IMB18_6200;
    -- flow-through select operator MUX_6647_inst
    IMC10_6648 <= IMB21_6224 when (BITSEL_u8_u1_6644_wire(0) /=  '0') else IMB20_6216;
    -- flow-through select operator MUX_6655_inst
    IMC11_6656 <= IMB23_6240 when (BITSEL_u8_u1_6652_wire(0) /=  '0') else IMB22_6232;
    -- flow-through select operator MUX_6663_inst
    IMC12_6664 <= IMB25_6256 when (BITSEL_u8_u1_6660_wire(0) /=  '0') else IMB24_6248;
    -- flow-through select operator MUX_6671_inst
    IMC13_6672 <= IMB27_6272 when (BITSEL_u8_u1_6668_wire(0) /=  '0') else IMB26_6264;
    -- flow-through select operator MUX_6679_inst
    IMC14_6680 <= IMB29_6288 when (BITSEL_u8_u1_6676_wire(0) /=  '0') else IMB28_6280;
    -- flow-through select operator MUX_6687_inst
    IMC15_6688 <= IMB31_6304 when (BITSEL_u8_u1_6684_wire(0) /=  '0') else IMB30_6296;
    -- flow-through select operator MUX_6695_inst
    IMC16_6696 <= IMB33_6320 when (BITSEL_u8_u1_6692_wire(0) /=  '0') else IMB32_6312;
    -- flow-through select operator MUX_6703_inst
    IMC17_6704 <= IMB35_6336 when (BITSEL_u8_u1_6700_wire(0) /=  '0') else IMB34_6328;
    -- flow-through select operator MUX_6711_inst
    IMC18_6712 <= IMB37_6352 when (BITSEL_u8_u1_6708_wire(0) /=  '0') else IMB36_6344;
    -- flow-through select operator MUX_6719_inst
    IMC19_6720 <= IMB39_6368 when (BITSEL_u8_u1_6716_wire(0) /=  '0') else IMB38_6360;
    -- flow-through select operator MUX_6727_inst
    IMC20_6728 <= IMB41_6384 when (BITSEL_u8_u1_6724_wire(0) /=  '0') else IMB40_6376;
    -- flow-through select operator MUX_6735_inst
    IMC21_6736 <= IMB43_6400 when (BITSEL_u8_u1_6732_wire(0) /=  '0') else IMB42_6392;
    -- flow-through select operator MUX_6743_inst
    IMC22_6744 <= IMB45_6416 when (BITSEL_u8_u1_6740_wire(0) /=  '0') else IMB44_6408;
    -- flow-through select operator MUX_6751_inst
    IMC23_6752 <= IMB47_6432 when (BITSEL_u8_u1_6748_wire(0) /=  '0') else IMB46_6424;
    -- flow-through select operator MUX_6759_inst
    IMC24_6760 <= IMB49_6448 when (BITSEL_u8_u1_6756_wire(0) /=  '0') else IMB48_6440;
    -- flow-through select operator MUX_6767_inst
    IMC25_6768 <= IMB51_6464 when (BITSEL_u8_u1_6764_wire(0) /=  '0') else IMB50_6456;
    -- flow-through select operator MUX_6775_inst
    IMC26_6776 <= IMB53_6480 when (BITSEL_u8_u1_6772_wire(0) /=  '0') else IMB52_6472;
    -- flow-through select operator MUX_6783_inst
    IMC27_6784 <= IMB55_6496 when (BITSEL_u8_u1_6780_wire(0) /=  '0') else IMB54_6488;
    -- flow-through select operator MUX_6791_inst
    IMC28_6792 <= IMB57_6512 when (BITSEL_u8_u1_6788_wire(0) /=  '0') else IMB56_6504;
    -- flow-through select operator MUX_6799_inst
    IMC29_6800 <= IMB59_6528 when (BITSEL_u8_u1_6796_wire(0) /=  '0') else IMB58_6520;
    -- flow-through select operator MUX_6807_inst
    IMC30_6808 <= IMB61_6544 when (BITSEL_u8_u1_6804_wire(0) /=  '0') else IMB60_6536;
    -- flow-through select operator MUX_6815_inst
    IMC31_6816 <= IMB63_6560 when (BITSEL_u8_u1_6812_wire(0) /=  '0') else IMB62_6552;
    -- flow-through select operator MUX_6823_inst
    IMD0_6824 <= IMC1_6576 when (BITSEL_u8_u1_6820_wire(0) /=  '0') else IMC0_6568;
    -- flow-through select operator MUX_6831_inst
    IMD1_6832 <= IMC3_6592 when (BITSEL_u8_u1_6828_wire(0) /=  '0') else IMC2_6584;
    -- flow-through select operator MUX_6839_inst
    IMD2_6840 <= IMC5_6608 when (BITSEL_u8_u1_6836_wire(0) /=  '0') else IMC4_6600;
    -- flow-through select operator MUX_6847_inst
    IMD3_6848 <= IMC7_6624 when (BITSEL_u8_u1_6844_wire(0) /=  '0') else IMC6_6616;
    -- flow-through select operator MUX_6855_inst
    IMD4_6856 <= IMC9_6640 when (BITSEL_u8_u1_6852_wire(0) /=  '0') else IMC8_6632;
    -- flow-through select operator MUX_6863_inst
    IMD5_6864 <= IMC11_6656 when (BITSEL_u8_u1_6860_wire(0) /=  '0') else IMC10_6648;
    -- flow-through select operator MUX_6871_inst
    IMD6_6872 <= IMC13_6672 when (BITSEL_u8_u1_6868_wire(0) /=  '0') else IMC12_6664;
    -- flow-through select operator MUX_6879_inst
    IMD7_6880 <= IMC15_6688 when (BITSEL_u8_u1_6876_wire(0) /=  '0') else IMC14_6680;
    -- flow-through select operator MUX_6887_inst
    IMD8_6888 <= IMC17_6704 when (BITSEL_u8_u1_6884_wire(0) /=  '0') else IMC16_6696;
    -- flow-through select operator MUX_6895_inst
    IMD9_6896 <= IMC19_6720 when (BITSEL_u8_u1_6892_wire(0) /=  '0') else IMC18_6712;
    -- flow-through select operator MUX_6903_inst
    IMD10_6904 <= IMC21_6736 when (BITSEL_u8_u1_6900_wire(0) /=  '0') else IMC20_6728;
    -- flow-through select operator MUX_6911_inst
    IMD11_6912 <= IMC23_6752 when (BITSEL_u8_u1_6908_wire(0) /=  '0') else IMC22_6744;
    -- flow-through select operator MUX_6919_inst
    IMD12_6920 <= IMC25_6768 when (BITSEL_u8_u1_6916_wire(0) /=  '0') else IMC24_6760;
    -- flow-through select operator MUX_6927_inst
    IMD13_6928 <= IMC27_6784 when (BITSEL_u8_u1_6924_wire(0) /=  '0') else IMC26_6776;
    -- flow-through select operator MUX_6935_inst
    IMD14_6936 <= IMC29_6800 when (BITSEL_u8_u1_6932_wire(0) /=  '0') else IMC28_6792;
    -- flow-through select operator MUX_6943_inst
    IMD15_6944 <= IMC31_6816 when (BITSEL_u8_u1_6940_wire(0) /=  '0') else IMC30_6808;
    -- flow-through select operator MUX_6951_inst
    IME0_6952 <= IMD1_6832 when (BITSEL_u8_u1_6948_wire(0) /=  '0') else IMD0_6824;
    -- flow-through select operator MUX_6959_inst
    IME1_6960 <= IMD3_6848 when (BITSEL_u8_u1_6956_wire(0) /=  '0') else IMD2_6840;
    -- flow-through select operator MUX_6967_inst
    IME2_6968 <= IMD5_6864 when (BITSEL_u8_u1_6964_wire(0) /=  '0') else IMD4_6856;
    -- flow-through select operator MUX_6975_inst
    IME3_6976 <= IMD7_6880 when (BITSEL_u8_u1_6972_wire(0) /=  '0') else IMD6_6872;
    -- flow-through select operator MUX_6983_inst
    IME4_6984 <= IMD9_6896 when (BITSEL_u8_u1_6980_wire(0) /=  '0') else IMD8_6888;
    -- flow-through select operator MUX_6991_inst
    IME5_6992 <= IMD11_6912 when (BITSEL_u8_u1_6988_wire(0) /=  '0') else IMD10_6904;
    -- flow-through select operator MUX_6999_inst
    IME6_7000 <= IMD13_6928 when (BITSEL_u8_u1_6996_wire(0) /=  '0') else IMD12_6920;
    -- flow-through select operator MUX_7007_inst
    IME7_7008 <= IMD15_6944 when (BITSEL_u8_u1_7004_wire(0) /=  '0') else IMD14_6936;
    -- flow-through select operator MUX_7015_inst
    IMF0_7016 <= IME1_6960 when (BITSEL_u8_u1_7012_wire(0) /=  '0') else IME0_6952;
    -- flow-through select operator MUX_7023_inst
    IMF1_7024 <= IME3_6976 when (BITSEL_u8_u1_7020_wire(0) /=  '0') else IME2_6968;
    -- flow-through select operator MUX_7031_inst
    IMF2_7032 <= IME5_6992 when (BITSEL_u8_u1_7028_wire(0) /=  '0') else IME4_6984;
    -- flow-through select operator MUX_7039_inst
    IMF3_7040 <= IME7_7008 when (BITSEL_u8_u1_7036_wire(0) /=  '0') else IME6_7000;
    -- flow-through select operator MUX_7047_inst
    IMG0_7048 <= IMF1_7024 when (BITSEL_u8_u1_7044_wire(0) /=  '0') else IMF0_7016;
    -- flow-through select operator MUX_7055_inst
    IMG1_7056 <= IMF3_7040 when (BITSEL_u8_u1_7052_wire(0) /=  '0') else IMF2_7032;
    -- flow-through select operator MUX_7063_inst
    s_out_buffer <= IMG1_7056 when (BITSEL_u8_u1_7060_wire(0) /=  '0') else IMG0_7048;
    -- binary operator BITSEL_u8_u1_4772_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4771_wire_constant, tmp_var);
      BITSEL_u8_u1_4772_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4782_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4781_wire_constant, tmp_var);
      BITSEL_u8_u1_4782_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4792_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4791_wire_constant, tmp_var);
      BITSEL_u8_u1_4792_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4802_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4801_wire_constant, tmp_var);
      BITSEL_u8_u1_4802_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4812_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4811_wire_constant, tmp_var);
      BITSEL_u8_u1_4812_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4822_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4821_wire_constant, tmp_var);
      BITSEL_u8_u1_4822_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4832_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4831_wire_constant, tmp_var);
      BITSEL_u8_u1_4832_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4842_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4841_wire_constant, tmp_var);
      BITSEL_u8_u1_4842_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4852_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4851_wire_constant, tmp_var);
      BITSEL_u8_u1_4852_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4862_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4861_wire_constant, tmp_var);
      BITSEL_u8_u1_4862_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4872_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4871_wire_constant, tmp_var);
      BITSEL_u8_u1_4872_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4882_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4881_wire_constant, tmp_var);
      BITSEL_u8_u1_4882_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4892_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4891_wire_constant, tmp_var);
      BITSEL_u8_u1_4892_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4902_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4901_wire_constant, tmp_var);
      BITSEL_u8_u1_4902_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4912_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4911_wire_constant, tmp_var);
      BITSEL_u8_u1_4912_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4922_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4921_wire_constant, tmp_var);
      BITSEL_u8_u1_4922_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4932_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4931_wire_constant, tmp_var);
      BITSEL_u8_u1_4932_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4942_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4941_wire_constant, tmp_var);
      BITSEL_u8_u1_4942_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4952_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4951_wire_constant, tmp_var);
      BITSEL_u8_u1_4952_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4962_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4961_wire_constant, tmp_var);
      BITSEL_u8_u1_4962_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4972_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4971_wire_constant, tmp_var);
      BITSEL_u8_u1_4972_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4982_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4981_wire_constant, tmp_var);
      BITSEL_u8_u1_4982_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_4992_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_4991_wire_constant, tmp_var);
      BITSEL_u8_u1_4992_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_5002_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5001_wire_constant, tmp_var);
      BITSEL_u8_u1_5002_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_5012_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5011_wire_constant, tmp_var);
      BITSEL_u8_u1_5012_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_5022_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5021_wire_constant, tmp_var);
      BITSEL_u8_u1_5022_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_5032_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5031_wire_constant, tmp_var);
      BITSEL_u8_u1_5032_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_5042_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5041_wire_constant, tmp_var);
      BITSEL_u8_u1_5042_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_5052_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5051_wire_constant, tmp_var);
      BITSEL_u8_u1_5052_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_5062_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5061_wire_constant, tmp_var);
      BITSEL_u8_u1_5062_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_5072_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5071_wire_constant, tmp_var);
      BITSEL_u8_u1_5072_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_5082_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5081_wire_constant, tmp_var);
      BITSEL_u8_u1_5082_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_5092_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5091_wire_constant, tmp_var);
      BITSEL_u8_u1_5092_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_5102_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5101_wire_constant, tmp_var);
      BITSEL_u8_u1_5102_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_5112_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5111_wire_constant, tmp_var);
      BITSEL_u8_u1_5112_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_5122_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5121_wire_constant, tmp_var);
      BITSEL_u8_u1_5122_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_5132_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5131_wire_constant, tmp_var);
      BITSEL_u8_u1_5132_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_5142_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5141_wire_constant, tmp_var);
      BITSEL_u8_u1_5142_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_5152_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5151_wire_constant, tmp_var);
      BITSEL_u8_u1_5152_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_5162_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5161_wire_constant, tmp_var);
      BITSEL_u8_u1_5162_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_5172_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5171_wire_constant, tmp_var);
      BITSEL_u8_u1_5172_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_5182_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5181_wire_constant, tmp_var);
      BITSEL_u8_u1_5182_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_5192_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5191_wire_constant, tmp_var);
      BITSEL_u8_u1_5192_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_5202_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5201_wire_constant, tmp_var);
      BITSEL_u8_u1_5202_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_5212_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5211_wire_constant, tmp_var);
      BITSEL_u8_u1_5212_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_5222_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5221_wire_constant, tmp_var);
      BITSEL_u8_u1_5222_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_5232_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5231_wire_constant, tmp_var);
      BITSEL_u8_u1_5232_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_5242_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5241_wire_constant, tmp_var);
      BITSEL_u8_u1_5242_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_5252_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5251_wire_constant, tmp_var);
      BITSEL_u8_u1_5252_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_5262_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5261_wire_constant, tmp_var);
      BITSEL_u8_u1_5262_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_5272_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5271_wire_constant, tmp_var);
      BITSEL_u8_u1_5272_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_5282_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5281_wire_constant, tmp_var);
      BITSEL_u8_u1_5282_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_5292_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5291_wire_constant, tmp_var);
      BITSEL_u8_u1_5292_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_5302_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5301_wire_constant, tmp_var);
      BITSEL_u8_u1_5302_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_5312_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5311_wire_constant, tmp_var);
      BITSEL_u8_u1_5312_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_5322_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5321_wire_constant, tmp_var);
      BITSEL_u8_u1_5322_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_5332_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5331_wire_constant, tmp_var);
      BITSEL_u8_u1_5332_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_5342_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5341_wire_constant, tmp_var);
      BITSEL_u8_u1_5342_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_5352_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5351_wire_constant, tmp_var);
      BITSEL_u8_u1_5352_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_5362_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5361_wire_constant, tmp_var);
      BITSEL_u8_u1_5362_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_5372_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5371_wire_constant, tmp_var);
      BITSEL_u8_u1_5372_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_5382_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5381_wire_constant, tmp_var);
      BITSEL_u8_u1_5382_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_5392_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5391_wire_constant, tmp_var);
      BITSEL_u8_u1_5392_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_5402_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5401_wire_constant, tmp_var);
      BITSEL_u8_u1_5402_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_5412_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5411_wire_constant, tmp_var);
      BITSEL_u8_u1_5412_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_5422_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5421_wire_constant, tmp_var);
      BITSEL_u8_u1_5422_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_5432_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5431_wire_constant, tmp_var);
      BITSEL_u8_u1_5432_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_5442_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5441_wire_constant, tmp_var);
      BITSEL_u8_u1_5442_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_5452_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5451_wire_constant, tmp_var);
      BITSEL_u8_u1_5452_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_5462_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5461_wire_constant, tmp_var);
      BITSEL_u8_u1_5462_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_5472_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5471_wire_constant, tmp_var);
      BITSEL_u8_u1_5472_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_5482_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5481_wire_constant, tmp_var);
      BITSEL_u8_u1_5482_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_5492_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5491_wire_constant, tmp_var);
      BITSEL_u8_u1_5492_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_5502_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5501_wire_constant, tmp_var);
      BITSEL_u8_u1_5502_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_5512_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5511_wire_constant, tmp_var);
      BITSEL_u8_u1_5512_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_5522_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5521_wire_constant, tmp_var);
      BITSEL_u8_u1_5522_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_5532_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5531_wire_constant, tmp_var);
      BITSEL_u8_u1_5532_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_5542_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5541_wire_constant, tmp_var);
      BITSEL_u8_u1_5542_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_5552_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5551_wire_constant, tmp_var);
      BITSEL_u8_u1_5552_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_5562_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5561_wire_constant, tmp_var);
      BITSEL_u8_u1_5562_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_5572_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5571_wire_constant, tmp_var);
      BITSEL_u8_u1_5572_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_5582_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5581_wire_constant, tmp_var);
      BITSEL_u8_u1_5582_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_5592_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5591_wire_constant, tmp_var);
      BITSEL_u8_u1_5592_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_5602_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5601_wire_constant, tmp_var);
      BITSEL_u8_u1_5602_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_5612_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5611_wire_constant, tmp_var);
      BITSEL_u8_u1_5612_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_5622_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5621_wire_constant, tmp_var);
      BITSEL_u8_u1_5622_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_5632_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5631_wire_constant, tmp_var);
      BITSEL_u8_u1_5632_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_5642_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5641_wire_constant, tmp_var);
      BITSEL_u8_u1_5642_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_5652_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5651_wire_constant, tmp_var);
      BITSEL_u8_u1_5652_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_5662_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5661_wire_constant, tmp_var);
      BITSEL_u8_u1_5662_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_5672_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5671_wire_constant, tmp_var);
      BITSEL_u8_u1_5672_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_5682_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5681_wire_constant, tmp_var);
      BITSEL_u8_u1_5682_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_5692_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5691_wire_constant, tmp_var);
      BITSEL_u8_u1_5692_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_5702_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5701_wire_constant, tmp_var);
      BITSEL_u8_u1_5702_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_5712_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5711_wire_constant, tmp_var);
      BITSEL_u8_u1_5712_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_5722_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5721_wire_constant, tmp_var);
      BITSEL_u8_u1_5722_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_5732_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5731_wire_constant, tmp_var);
      BITSEL_u8_u1_5732_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_5742_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5741_wire_constant, tmp_var);
      BITSEL_u8_u1_5742_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_5752_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5751_wire_constant, tmp_var);
      BITSEL_u8_u1_5752_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_5762_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5761_wire_constant, tmp_var);
      BITSEL_u8_u1_5762_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_5772_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5771_wire_constant, tmp_var);
      BITSEL_u8_u1_5772_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_5782_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5781_wire_constant, tmp_var);
      BITSEL_u8_u1_5782_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_5792_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5791_wire_constant, tmp_var);
      BITSEL_u8_u1_5792_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_5802_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5801_wire_constant, tmp_var);
      BITSEL_u8_u1_5802_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_5812_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5811_wire_constant, tmp_var);
      BITSEL_u8_u1_5812_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_5822_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5821_wire_constant, tmp_var);
      BITSEL_u8_u1_5822_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_5832_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5831_wire_constant, tmp_var);
      BITSEL_u8_u1_5832_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_5842_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5841_wire_constant, tmp_var);
      BITSEL_u8_u1_5842_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_5852_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5851_wire_constant, tmp_var);
      BITSEL_u8_u1_5852_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_5862_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5861_wire_constant, tmp_var);
      BITSEL_u8_u1_5862_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_5872_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5871_wire_constant, tmp_var);
      BITSEL_u8_u1_5872_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_5882_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5881_wire_constant, tmp_var);
      BITSEL_u8_u1_5882_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_5892_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5891_wire_constant, tmp_var);
      BITSEL_u8_u1_5892_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_5902_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5901_wire_constant, tmp_var);
      BITSEL_u8_u1_5902_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_5912_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5911_wire_constant, tmp_var);
      BITSEL_u8_u1_5912_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_5922_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5921_wire_constant, tmp_var);
      BITSEL_u8_u1_5922_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_5932_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5931_wire_constant, tmp_var);
      BITSEL_u8_u1_5932_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_5942_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5941_wire_constant, tmp_var);
      BITSEL_u8_u1_5942_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_5952_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5951_wire_constant, tmp_var);
      BITSEL_u8_u1_5952_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_5962_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5961_wire_constant, tmp_var);
      BITSEL_u8_u1_5962_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_5972_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5971_wire_constant, tmp_var);
      BITSEL_u8_u1_5972_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_5982_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5981_wire_constant, tmp_var);
      BITSEL_u8_u1_5982_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_5992_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_5991_wire_constant, tmp_var);
      BITSEL_u8_u1_5992_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6002_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6001_wire_constant, tmp_var);
      BITSEL_u8_u1_6002_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6012_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6011_wire_constant, tmp_var);
      BITSEL_u8_u1_6012_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6022_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6021_wire_constant, tmp_var);
      BITSEL_u8_u1_6022_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6032_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6031_wire_constant, tmp_var);
      BITSEL_u8_u1_6032_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6042_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6041_wire_constant, tmp_var);
      BITSEL_u8_u1_6042_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6052_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6051_wire_constant, tmp_var);
      BITSEL_u8_u1_6052_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6060_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6059_wire_constant, tmp_var);
      BITSEL_u8_u1_6060_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6068_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6067_wire_constant, tmp_var);
      BITSEL_u8_u1_6068_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6076_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6075_wire_constant, tmp_var);
      BITSEL_u8_u1_6076_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6084_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6083_wire_constant, tmp_var);
      BITSEL_u8_u1_6084_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6092_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6091_wire_constant, tmp_var);
      BITSEL_u8_u1_6092_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6100_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6099_wire_constant, tmp_var);
      BITSEL_u8_u1_6100_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6108_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6107_wire_constant, tmp_var);
      BITSEL_u8_u1_6108_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6116_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6115_wire_constant, tmp_var);
      BITSEL_u8_u1_6116_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6124_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6123_wire_constant, tmp_var);
      BITSEL_u8_u1_6124_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6132_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6131_wire_constant, tmp_var);
      BITSEL_u8_u1_6132_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6140_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6139_wire_constant, tmp_var);
      BITSEL_u8_u1_6140_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6148_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6147_wire_constant, tmp_var);
      BITSEL_u8_u1_6148_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6156_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6155_wire_constant, tmp_var);
      BITSEL_u8_u1_6156_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6164_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6163_wire_constant, tmp_var);
      BITSEL_u8_u1_6164_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6172_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6171_wire_constant, tmp_var);
      BITSEL_u8_u1_6172_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6180_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6179_wire_constant, tmp_var);
      BITSEL_u8_u1_6180_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6188_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6187_wire_constant, tmp_var);
      BITSEL_u8_u1_6188_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6196_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6195_wire_constant, tmp_var);
      BITSEL_u8_u1_6196_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6204_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6203_wire_constant, tmp_var);
      BITSEL_u8_u1_6204_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6212_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6211_wire_constant, tmp_var);
      BITSEL_u8_u1_6212_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6220_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6219_wire_constant, tmp_var);
      BITSEL_u8_u1_6220_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6228_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6227_wire_constant, tmp_var);
      BITSEL_u8_u1_6228_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6236_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6235_wire_constant, tmp_var);
      BITSEL_u8_u1_6236_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6244_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6243_wire_constant, tmp_var);
      BITSEL_u8_u1_6244_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6252_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6251_wire_constant, tmp_var);
      BITSEL_u8_u1_6252_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6260_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6259_wire_constant, tmp_var);
      BITSEL_u8_u1_6260_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6268_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6267_wire_constant, tmp_var);
      BITSEL_u8_u1_6268_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6276_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6275_wire_constant, tmp_var);
      BITSEL_u8_u1_6276_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6284_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6283_wire_constant, tmp_var);
      BITSEL_u8_u1_6284_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6292_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6291_wire_constant, tmp_var);
      BITSEL_u8_u1_6292_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6300_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6299_wire_constant, tmp_var);
      BITSEL_u8_u1_6300_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6308_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6307_wire_constant, tmp_var);
      BITSEL_u8_u1_6308_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6316_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6315_wire_constant, tmp_var);
      BITSEL_u8_u1_6316_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6324_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6323_wire_constant, tmp_var);
      BITSEL_u8_u1_6324_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6332_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6331_wire_constant, tmp_var);
      BITSEL_u8_u1_6332_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6340_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6339_wire_constant, tmp_var);
      BITSEL_u8_u1_6340_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6348_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6347_wire_constant, tmp_var);
      BITSEL_u8_u1_6348_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6356_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6355_wire_constant, tmp_var);
      BITSEL_u8_u1_6356_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6364_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6363_wire_constant, tmp_var);
      BITSEL_u8_u1_6364_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6372_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6371_wire_constant, tmp_var);
      BITSEL_u8_u1_6372_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6380_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6379_wire_constant, tmp_var);
      BITSEL_u8_u1_6380_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6388_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6387_wire_constant, tmp_var);
      BITSEL_u8_u1_6388_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6396_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6395_wire_constant, tmp_var);
      BITSEL_u8_u1_6396_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6404_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6403_wire_constant, tmp_var);
      BITSEL_u8_u1_6404_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6412_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6411_wire_constant, tmp_var);
      BITSEL_u8_u1_6412_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6420_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6419_wire_constant, tmp_var);
      BITSEL_u8_u1_6420_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6428_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6427_wire_constant, tmp_var);
      BITSEL_u8_u1_6428_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6436_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6435_wire_constant, tmp_var);
      BITSEL_u8_u1_6436_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6444_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6443_wire_constant, tmp_var);
      BITSEL_u8_u1_6444_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6452_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6451_wire_constant, tmp_var);
      BITSEL_u8_u1_6452_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6460_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6459_wire_constant, tmp_var);
      BITSEL_u8_u1_6460_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6468_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6467_wire_constant, tmp_var);
      BITSEL_u8_u1_6468_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6476_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6475_wire_constant, tmp_var);
      BITSEL_u8_u1_6476_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6484_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6483_wire_constant, tmp_var);
      BITSEL_u8_u1_6484_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6492_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6491_wire_constant, tmp_var);
      BITSEL_u8_u1_6492_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6500_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6499_wire_constant, tmp_var);
      BITSEL_u8_u1_6500_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6508_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6507_wire_constant, tmp_var);
      BITSEL_u8_u1_6508_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6516_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6515_wire_constant, tmp_var);
      BITSEL_u8_u1_6516_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6524_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6523_wire_constant, tmp_var);
      BITSEL_u8_u1_6524_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6532_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6531_wire_constant, tmp_var);
      BITSEL_u8_u1_6532_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6540_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6539_wire_constant, tmp_var);
      BITSEL_u8_u1_6540_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6548_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6547_wire_constant, tmp_var);
      BITSEL_u8_u1_6548_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6556_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6555_wire_constant, tmp_var);
      BITSEL_u8_u1_6556_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6564_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6563_wire_constant, tmp_var);
      BITSEL_u8_u1_6564_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6572_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6571_wire_constant, tmp_var);
      BITSEL_u8_u1_6572_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6580_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6579_wire_constant, tmp_var);
      BITSEL_u8_u1_6580_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6588_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6587_wire_constant, tmp_var);
      BITSEL_u8_u1_6588_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6596_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6595_wire_constant, tmp_var);
      BITSEL_u8_u1_6596_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6604_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6603_wire_constant, tmp_var);
      BITSEL_u8_u1_6604_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6612_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6611_wire_constant, tmp_var);
      BITSEL_u8_u1_6612_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6620_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6619_wire_constant, tmp_var);
      BITSEL_u8_u1_6620_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6628_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6627_wire_constant, tmp_var);
      BITSEL_u8_u1_6628_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6636_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6635_wire_constant, tmp_var);
      BITSEL_u8_u1_6636_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6644_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6643_wire_constant, tmp_var);
      BITSEL_u8_u1_6644_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6652_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6651_wire_constant, tmp_var);
      BITSEL_u8_u1_6652_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6660_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6659_wire_constant, tmp_var);
      BITSEL_u8_u1_6660_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6668_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6667_wire_constant, tmp_var);
      BITSEL_u8_u1_6668_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6676_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6675_wire_constant, tmp_var);
      BITSEL_u8_u1_6676_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6684_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6683_wire_constant, tmp_var);
      BITSEL_u8_u1_6684_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6692_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6691_wire_constant, tmp_var);
      BITSEL_u8_u1_6692_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6700_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6699_wire_constant, tmp_var);
      BITSEL_u8_u1_6700_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6708_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6707_wire_constant, tmp_var);
      BITSEL_u8_u1_6708_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6716_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6715_wire_constant, tmp_var);
      BITSEL_u8_u1_6716_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6724_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6723_wire_constant, tmp_var);
      BITSEL_u8_u1_6724_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6732_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6731_wire_constant, tmp_var);
      BITSEL_u8_u1_6732_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6740_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6739_wire_constant, tmp_var);
      BITSEL_u8_u1_6740_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6748_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6747_wire_constant, tmp_var);
      BITSEL_u8_u1_6748_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6756_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6755_wire_constant, tmp_var);
      BITSEL_u8_u1_6756_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6764_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6763_wire_constant, tmp_var);
      BITSEL_u8_u1_6764_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6772_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6771_wire_constant, tmp_var);
      BITSEL_u8_u1_6772_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6780_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6779_wire_constant, tmp_var);
      BITSEL_u8_u1_6780_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6788_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6787_wire_constant, tmp_var);
      BITSEL_u8_u1_6788_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6796_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6795_wire_constant, tmp_var);
      BITSEL_u8_u1_6796_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6804_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6803_wire_constant, tmp_var);
      BITSEL_u8_u1_6804_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6812_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6811_wire_constant, tmp_var);
      BITSEL_u8_u1_6812_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6820_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6819_wire_constant, tmp_var);
      BITSEL_u8_u1_6820_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6828_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6827_wire_constant, tmp_var);
      BITSEL_u8_u1_6828_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6836_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6835_wire_constant, tmp_var);
      BITSEL_u8_u1_6836_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6844_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6843_wire_constant, tmp_var);
      BITSEL_u8_u1_6844_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6852_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6851_wire_constant, tmp_var);
      BITSEL_u8_u1_6852_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6860_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6859_wire_constant, tmp_var);
      BITSEL_u8_u1_6860_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6868_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6867_wire_constant, tmp_var);
      BITSEL_u8_u1_6868_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6876_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6875_wire_constant, tmp_var);
      BITSEL_u8_u1_6876_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6884_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6883_wire_constant, tmp_var);
      BITSEL_u8_u1_6884_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6892_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6891_wire_constant, tmp_var);
      BITSEL_u8_u1_6892_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6900_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6899_wire_constant, tmp_var);
      BITSEL_u8_u1_6900_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6908_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6907_wire_constant, tmp_var);
      BITSEL_u8_u1_6908_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6916_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6915_wire_constant, tmp_var);
      BITSEL_u8_u1_6916_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6924_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6923_wire_constant, tmp_var);
      BITSEL_u8_u1_6924_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6932_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6931_wire_constant, tmp_var);
      BITSEL_u8_u1_6932_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6940_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6939_wire_constant, tmp_var);
      BITSEL_u8_u1_6940_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6948_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6947_wire_constant, tmp_var);
      BITSEL_u8_u1_6948_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6956_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6955_wire_constant, tmp_var);
      BITSEL_u8_u1_6956_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6964_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6963_wire_constant, tmp_var);
      BITSEL_u8_u1_6964_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6972_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6971_wire_constant, tmp_var);
      BITSEL_u8_u1_6972_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6980_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6979_wire_constant, tmp_var);
      BITSEL_u8_u1_6980_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6988_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6987_wire_constant, tmp_var);
      BITSEL_u8_u1_6988_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_6996_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_6995_wire_constant, tmp_var);
      BITSEL_u8_u1_6996_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_7004_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7003_wire_constant, tmp_var);
      BITSEL_u8_u1_7004_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_7012_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7011_wire_constant, tmp_var);
      BITSEL_u8_u1_7012_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_7020_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7019_wire_constant, tmp_var);
      BITSEL_u8_u1_7020_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_7028_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7027_wire_constant, tmp_var);
      BITSEL_u8_u1_7028_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_7036_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7035_wire_constant, tmp_var);
      BITSEL_u8_u1_7036_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_7044_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7043_wire_constant, tmp_var);
      BITSEL_u8_u1_7044_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_7052_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7051_wire_constant, tmp_var);
      BITSEL_u8_u1_7052_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_7060_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7059_wire_constant, tmp_var);
      BITSEL_u8_u1_7060_wire <= tmp_var; -- 
    end process;
    -- 
  end Block; -- data_path
  -- 
end Inv_Sbox_3_Volatile_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library work;
use work.ahir_system_global_package.all;
entity Inv_Sbox_4_Volatile is -- 
  port ( -- 
    s_in : in  std_logic_vector(7 downto 0);
    s_out : out  std_logic_vector(7 downto 0)-- 
  );
  -- 
end entity Inv_Sbox_4_Volatile;
architecture Inv_Sbox_4_Volatile_arch of Inv_Sbox_4_Volatile is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector(8-1 downto 0);
  signal default_zero_sig: std_logic;
  -- input port buffer signals
  signal s_in_buffer :  std_logic_vector(7 downto 0);
  -- output port buffer signals
  signal s_out_buffer :  std_logic_vector(7 downto 0);
  -- volatile/operator module components. 
  -- 
begin --  
  -- input handling ------------------------------------------------
  s_in_buffer <= s_in;
  -- output handling  -------------------------------------------------------
  s_out <= s_out_buffer;
  -- the control path --------------------------------------------------
  default_zero_sig <= '0';
  -- volatile module, no control path
  -- the data path
  data_path: Block -- 
    signal BITSEL_u8_u1_7072_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7082_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7092_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7102_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7112_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7122_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7132_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7142_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7152_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7162_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7172_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7182_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7192_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7202_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7212_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7222_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7232_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7242_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7252_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7262_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7272_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7282_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7292_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7302_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7312_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7322_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7332_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7342_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7352_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7362_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7372_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7382_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7392_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7402_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7412_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7422_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7432_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7442_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7452_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7462_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7472_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7482_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7492_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7502_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7512_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7522_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7532_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7542_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7552_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7562_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7572_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7582_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7592_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7602_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7612_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7622_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7632_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7642_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7652_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7662_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7672_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7682_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7692_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7702_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7712_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7722_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7732_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7742_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7752_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7762_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7772_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7782_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7792_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7802_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7812_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7822_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7832_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7842_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7852_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7862_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7872_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7882_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7892_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7902_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7912_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7922_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7932_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7942_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7952_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7962_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7972_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7982_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_7992_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8002_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8012_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8022_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8032_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8042_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8052_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8062_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8072_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8082_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8092_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8102_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8112_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8122_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8132_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8142_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8152_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8162_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8172_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8182_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8192_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8202_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8212_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8222_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8232_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8242_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8252_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8262_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8272_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8282_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8292_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8302_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8312_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8322_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8332_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8342_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8352_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8360_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8368_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8376_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8384_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8392_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8400_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8408_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8416_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8424_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8432_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8440_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8448_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8456_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8464_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8472_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8480_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8488_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8496_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8504_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8512_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8520_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8528_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8536_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8544_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8552_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8560_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8568_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8576_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8584_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8592_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8600_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8608_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8616_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8624_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8632_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8640_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8648_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8656_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8664_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8672_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8680_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8688_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8696_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8704_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8712_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8720_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8728_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8736_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8744_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8752_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8760_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8768_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8776_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8784_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8792_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8800_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8808_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8816_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8824_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8832_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8840_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8848_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8856_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8864_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8872_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8880_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8888_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8896_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8904_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8912_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8920_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8928_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8936_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8944_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8952_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8960_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8968_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8976_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8984_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_8992_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9000_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9008_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9016_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9024_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9032_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9040_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9048_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9056_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9064_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9072_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9080_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9088_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9096_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9104_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9112_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9120_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9128_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9136_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9144_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9152_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9160_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9168_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9176_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9184_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9192_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9200_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9208_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9216_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9224_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9232_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9240_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9248_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9256_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9264_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9272_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9280_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9288_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9296_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9304_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9312_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9320_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9328_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9336_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9344_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9352_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9360_wire : std_logic_vector(0 downto 0);
    signal IMA0_7078 : std_logic_vector(7 downto 0);
    signal IMA100_8078 : std_logic_vector(7 downto 0);
    signal IMA101_8088 : std_logic_vector(7 downto 0);
    signal IMA102_8098 : std_logic_vector(7 downto 0);
    signal IMA103_8108 : std_logic_vector(7 downto 0);
    signal IMA104_8118 : std_logic_vector(7 downto 0);
    signal IMA105_8128 : std_logic_vector(7 downto 0);
    signal IMA106_8138 : std_logic_vector(7 downto 0);
    signal IMA107_8148 : std_logic_vector(7 downto 0);
    signal IMA108_8158 : std_logic_vector(7 downto 0);
    signal IMA109_8168 : std_logic_vector(7 downto 0);
    signal IMA10_7178 : std_logic_vector(7 downto 0);
    signal IMA110_8178 : std_logic_vector(7 downto 0);
    signal IMA111_8188 : std_logic_vector(7 downto 0);
    signal IMA112_8198 : std_logic_vector(7 downto 0);
    signal IMA113_8208 : std_logic_vector(7 downto 0);
    signal IMA114_8218 : std_logic_vector(7 downto 0);
    signal IMA115_8228 : std_logic_vector(7 downto 0);
    signal IMA116_8238 : std_logic_vector(7 downto 0);
    signal IMA117_8248 : std_logic_vector(7 downto 0);
    signal IMA118_8258 : std_logic_vector(7 downto 0);
    signal IMA119_8268 : std_logic_vector(7 downto 0);
    signal IMA11_7188 : std_logic_vector(7 downto 0);
    signal IMA120_8278 : std_logic_vector(7 downto 0);
    signal IMA121_8288 : std_logic_vector(7 downto 0);
    signal IMA122_8298 : std_logic_vector(7 downto 0);
    signal IMA123_8308 : std_logic_vector(7 downto 0);
    signal IMA124_8318 : std_logic_vector(7 downto 0);
    signal IMA125_8328 : std_logic_vector(7 downto 0);
    signal IMA126_8338 : std_logic_vector(7 downto 0);
    signal IMA127_8348 : std_logic_vector(7 downto 0);
    signal IMA12_7198 : std_logic_vector(7 downto 0);
    signal IMA13_7208 : std_logic_vector(7 downto 0);
    signal IMA14_7218 : std_logic_vector(7 downto 0);
    signal IMA15_7228 : std_logic_vector(7 downto 0);
    signal IMA16_7238 : std_logic_vector(7 downto 0);
    signal IMA17_7248 : std_logic_vector(7 downto 0);
    signal IMA18_7258 : std_logic_vector(7 downto 0);
    signal IMA19_7268 : std_logic_vector(7 downto 0);
    signal IMA1_7088 : std_logic_vector(7 downto 0);
    signal IMA20_7278 : std_logic_vector(7 downto 0);
    signal IMA21_7288 : std_logic_vector(7 downto 0);
    signal IMA22_7298 : std_logic_vector(7 downto 0);
    signal IMA23_7308 : std_logic_vector(7 downto 0);
    signal IMA24_7318 : std_logic_vector(7 downto 0);
    signal IMA25_7328 : std_logic_vector(7 downto 0);
    signal IMA26_7338 : std_logic_vector(7 downto 0);
    signal IMA27_7348 : std_logic_vector(7 downto 0);
    signal IMA28_7358 : std_logic_vector(7 downto 0);
    signal IMA29_7368 : std_logic_vector(7 downto 0);
    signal IMA2_7098 : std_logic_vector(7 downto 0);
    signal IMA30_7378 : std_logic_vector(7 downto 0);
    signal IMA31_7388 : std_logic_vector(7 downto 0);
    signal IMA32_7398 : std_logic_vector(7 downto 0);
    signal IMA33_7408 : std_logic_vector(7 downto 0);
    signal IMA34_7418 : std_logic_vector(7 downto 0);
    signal IMA35_7428 : std_logic_vector(7 downto 0);
    signal IMA36_7438 : std_logic_vector(7 downto 0);
    signal IMA37_7448 : std_logic_vector(7 downto 0);
    signal IMA38_7458 : std_logic_vector(7 downto 0);
    signal IMA39_7468 : std_logic_vector(7 downto 0);
    signal IMA3_7108 : std_logic_vector(7 downto 0);
    signal IMA40_7478 : std_logic_vector(7 downto 0);
    signal IMA41_7488 : std_logic_vector(7 downto 0);
    signal IMA42_7498 : std_logic_vector(7 downto 0);
    signal IMA43_7508 : std_logic_vector(7 downto 0);
    signal IMA44_7518 : std_logic_vector(7 downto 0);
    signal IMA45_7528 : std_logic_vector(7 downto 0);
    signal IMA46_7538 : std_logic_vector(7 downto 0);
    signal IMA47_7548 : std_logic_vector(7 downto 0);
    signal IMA48_7558 : std_logic_vector(7 downto 0);
    signal IMA49_7568 : std_logic_vector(7 downto 0);
    signal IMA4_7118 : std_logic_vector(7 downto 0);
    signal IMA50_7578 : std_logic_vector(7 downto 0);
    signal IMA51_7588 : std_logic_vector(7 downto 0);
    signal IMA52_7598 : std_logic_vector(7 downto 0);
    signal IMA53_7608 : std_logic_vector(7 downto 0);
    signal IMA54_7618 : std_logic_vector(7 downto 0);
    signal IMA55_7628 : std_logic_vector(7 downto 0);
    signal IMA56_7638 : std_logic_vector(7 downto 0);
    signal IMA57_7648 : std_logic_vector(7 downto 0);
    signal IMA58_7658 : std_logic_vector(7 downto 0);
    signal IMA59_7668 : std_logic_vector(7 downto 0);
    signal IMA5_7128 : std_logic_vector(7 downto 0);
    signal IMA60_7678 : std_logic_vector(7 downto 0);
    signal IMA61_7688 : std_logic_vector(7 downto 0);
    signal IMA62_7698 : std_logic_vector(7 downto 0);
    signal IMA63_7708 : std_logic_vector(7 downto 0);
    signal IMA64_7718 : std_logic_vector(7 downto 0);
    signal IMA65_7728 : std_logic_vector(7 downto 0);
    signal IMA66_7738 : std_logic_vector(7 downto 0);
    signal IMA67_7748 : std_logic_vector(7 downto 0);
    signal IMA68_7758 : std_logic_vector(7 downto 0);
    signal IMA69_7768 : std_logic_vector(7 downto 0);
    signal IMA6_7138 : std_logic_vector(7 downto 0);
    signal IMA70_7778 : std_logic_vector(7 downto 0);
    signal IMA71_7788 : std_logic_vector(7 downto 0);
    signal IMA72_7798 : std_logic_vector(7 downto 0);
    signal IMA73_7808 : std_logic_vector(7 downto 0);
    signal IMA74_7818 : std_logic_vector(7 downto 0);
    signal IMA75_7828 : std_logic_vector(7 downto 0);
    signal IMA76_7838 : std_logic_vector(7 downto 0);
    signal IMA77_7848 : std_logic_vector(7 downto 0);
    signal IMA78_7858 : std_logic_vector(7 downto 0);
    signal IMA79_7868 : std_logic_vector(7 downto 0);
    signal IMA7_7148 : std_logic_vector(7 downto 0);
    signal IMA80_7878 : std_logic_vector(7 downto 0);
    signal IMA81_7888 : std_logic_vector(7 downto 0);
    signal IMA82_7898 : std_logic_vector(7 downto 0);
    signal IMA83_7908 : std_logic_vector(7 downto 0);
    signal IMA84_7918 : std_logic_vector(7 downto 0);
    signal IMA85_7928 : std_logic_vector(7 downto 0);
    signal IMA86_7938 : std_logic_vector(7 downto 0);
    signal IMA87_7948 : std_logic_vector(7 downto 0);
    signal IMA88_7958 : std_logic_vector(7 downto 0);
    signal IMA89_7968 : std_logic_vector(7 downto 0);
    signal IMA8_7158 : std_logic_vector(7 downto 0);
    signal IMA90_7978 : std_logic_vector(7 downto 0);
    signal IMA91_7988 : std_logic_vector(7 downto 0);
    signal IMA92_7998 : std_logic_vector(7 downto 0);
    signal IMA93_8008 : std_logic_vector(7 downto 0);
    signal IMA94_8018 : std_logic_vector(7 downto 0);
    signal IMA95_8028 : std_logic_vector(7 downto 0);
    signal IMA96_8038 : std_logic_vector(7 downto 0);
    signal IMA97_8048 : std_logic_vector(7 downto 0);
    signal IMA98_8058 : std_logic_vector(7 downto 0);
    signal IMA99_8068 : std_logic_vector(7 downto 0);
    signal IMA9_7168 : std_logic_vector(7 downto 0);
    signal IMB0_8356 : std_logic_vector(7 downto 0);
    signal IMB10_8436 : std_logic_vector(7 downto 0);
    signal IMB11_8444 : std_logic_vector(7 downto 0);
    signal IMB12_8452 : std_logic_vector(7 downto 0);
    signal IMB13_8460 : std_logic_vector(7 downto 0);
    signal IMB14_8468 : std_logic_vector(7 downto 0);
    signal IMB15_8476 : std_logic_vector(7 downto 0);
    signal IMB16_8484 : std_logic_vector(7 downto 0);
    signal IMB17_8492 : std_logic_vector(7 downto 0);
    signal IMB18_8500 : std_logic_vector(7 downto 0);
    signal IMB19_8508 : std_logic_vector(7 downto 0);
    signal IMB1_8364 : std_logic_vector(7 downto 0);
    signal IMB20_8516 : std_logic_vector(7 downto 0);
    signal IMB21_8524 : std_logic_vector(7 downto 0);
    signal IMB22_8532 : std_logic_vector(7 downto 0);
    signal IMB23_8540 : std_logic_vector(7 downto 0);
    signal IMB24_8548 : std_logic_vector(7 downto 0);
    signal IMB25_8556 : std_logic_vector(7 downto 0);
    signal IMB26_8564 : std_logic_vector(7 downto 0);
    signal IMB27_8572 : std_logic_vector(7 downto 0);
    signal IMB28_8580 : std_logic_vector(7 downto 0);
    signal IMB29_8588 : std_logic_vector(7 downto 0);
    signal IMB2_8372 : std_logic_vector(7 downto 0);
    signal IMB30_8596 : std_logic_vector(7 downto 0);
    signal IMB31_8604 : std_logic_vector(7 downto 0);
    signal IMB32_8612 : std_logic_vector(7 downto 0);
    signal IMB33_8620 : std_logic_vector(7 downto 0);
    signal IMB34_8628 : std_logic_vector(7 downto 0);
    signal IMB35_8636 : std_logic_vector(7 downto 0);
    signal IMB36_8644 : std_logic_vector(7 downto 0);
    signal IMB37_8652 : std_logic_vector(7 downto 0);
    signal IMB38_8660 : std_logic_vector(7 downto 0);
    signal IMB39_8668 : std_logic_vector(7 downto 0);
    signal IMB3_8380 : std_logic_vector(7 downto 0);
    signal IMB40_8676 : std_logic_vector(7 downto 0);
    signal IMB41_8684 : std_logic_vector(7 downto 0);
    signal IMB42_8692 : std_logic_vector(7 downto 0);
    signal IMB43_8700 : std_logic_vector(7 downto 0);
    signal IMB44_8708 : std_logic_vector(7 downto 0);
    signal IMB45_8716 : std_logic_vector(7 downto 0);
    signal IMB46_8724 : std_logic_vector(7 downto 0);
    signal IMB47_8732 : std_logic_vector(7 downto 0);
    signal IMB48_8740 : std_logic_vector(7 downto 0);
    signal IMB49_8748 : std_logic_vector(7 downto 0);
    signal IMB4_8388 : std_logic_vector(7 downto 0);
    signal IMB50_8756 : std_logic_vector(7 downto 0);
    signal IMB51_8764 : std_logic_vector(7 downto 0);
    signal IMB52_8772 : std_logic_vector(7 downto 0);
    signal IMB53_8780 : std_logic_vector(7 downto 0);
    signal IMB54_8788 : std_logic_vector(7 downto 0);
    signal IMB55_8796 : std_logic_vector(7 downto 0);
    signal IMB56_8804 : std_logic_vector(7 downto 0);
    signal IMB57_8812 : std_logic_vector(7 downto 0);
    signal IMB58_8820 : std_logic_vector(7 downto 0);
    signal IMB59_8828 : std_logic_vector(7 downto 0);
    signal IMB5_8396 : std_logic_vector(7 downto 0);
    signal IMB60_8836 : std_logic_vector(7 downto 0);
    signal IMB61_8844 : std_logic_vector(7 downto 0);
    signal IMB62_8852 : std_logic_vector(7 downto 0);
    signal IMB63_8860 : std_logic_vector(7 downto 0);
    signal IMB6_8404 : std_logic_vector(7 downto 0);
    signal IMB7_8412 : std_logic_vector(7 downto 0);
    signal IMB8_8420 : std_logic_vector(7 downto 0);
    signal IMB9_8428 : std_logic_vector(7 downto 0);
    signal IMC0_8868 : std_logic_vector(7 downto 0);
    signal IMC10_8948 : std_logic_vector(7 downto 0);
    signal IMC11_8956 : std_logic_vector(7 downto 0);
    signal IMC12_8964 : std_logic_vector(7 downto 0);
    signal IMC13_8972 : std_logic_vector(7 downto 0);
    signal IMC14_8980 : std_logic_vector(7 downto 0);
    signal IMC15_8988 : std_logic_vector(7 downto 0);
    signal IMC16_8996 : std_logic_vector(7 downto 0);
    signal IMC17_9004 : std_logic_vector(7 downto 0);
    signal IMC18_9012 : std_logic_vector(7 downto 0);
    signal IMC19_9020 : std_logic_vector(7 downto 0);
    signal IMC1_8876 : std_logic_vector(7 downto 0);
    signal IMC20_9028 : std_logic_vector(7 downto 0);
    signal IMC21_9036 : std_logic_vector(7 downto 0);
    signal IMC22_9044 : std_logic_vector(7 downto 0);
    signal IMC23_9052 : std_logic_vector(7 downto 0);
    signal IMC24_9060 : std_logic_vector(7 downto 0);
    signal IMC25_9068 : std_logic_vector(7 downto 0);
    signal IMC26_9076 : std_logic_vector(7 downto 0);
    signal IMC27_9084 : std_logic_vector(7 downto 0);
    signal IMC28_9092 : std_logic_vector(7 downto 0);
    signal IMC29_9100 : std_logic_vector(7 downto 0);
    signal IMC2_8884 : std_logic_vector(7 downto 0);
    signal IMC30_9108 : std_logic_vector(7 downto 0);
    signal IMC31_9116 : std_logic_vector(7 downto 0);
    signal IMC3_8892 : std_logic_vector(7 downto 0);
    signal IMC4_8900 : std_logic_vector(7 downto 0);
    signal IMC5_8908 : std_logic_vector(7 downto 0);
    signal IMC6_8916 : std_logic_vector(7 downto 0);
    signal IMC7_8924 : std_logic_vector(7 downto 0);
    signal IMC8_8932 : std_logic_vector(7 downto 0);
    signal IMC9_8940 : std_logic_vector(7 downto 0);
    signal IMD0_9124 : std_logic_vector(7 downto 0);
    signal IMD10_9204 : std_logic_vector(7 downto 0);
    signal IMD11_9212 : std_logic_vector(7 downto 0);
    signal IMD12_9220 : std_logic_vector(7 downto 0);
    signal IMD13_9228 : std_logic_vector(7 downto 0);
    signal IMD14_9236 : std_logic_vector(7 downto 0);
    signal IMD15_9244 : std_logic_vector(7 downto 0);
    signal IMD1_9132 : std_logic_vector(7 downto 0);
    signal IMD2_9140 : std_logic_vector(7 downto 0);
    signal IMD3_9148 : std_logic_vector(7 downto 0);
    signal IMD4_9156 : std_logic_vector(7 downto 0);
    signal IMD5_9164 : std_logic_vector(7 downto 0);
    signal IMD6_9172 : std_logic_vector(7 downto 0);
    signal IMD7_9180 : std_logic_vector(7 downto 0);
    signal IMD8_9188 : std_logic_vector(7 downto 0);
    signal IMD9_9196 : std_logic_vector(7 downto 0);
    signal IME0_9252 : std_logic_vector(7 downto 0);
    signal IME1_9260 : std_logic_vector(7 downto 0);
    signal IME2_9268 : std_logic_vector(7 downto 0);
    signal IME3_9276 : std_logic_vector(7 downto 0);
    signal IME4_9284 : std_logic_vector(7 downto 0);
    signal IME5_9292 : std_logic_vector(7 downto 0);
    signal IME6_9300 : std_logic_vector(7 downto 0);
    signal IME7_9308 : std_logic_vector(7 downto 0);
    signal IMF0_9316 : std_logic_vector(7 downto 0);
    signal IMF1_9324 : std_logic_vector(7 downto 0);
    signal IMF2_9332 : std_logic_vector(7 downto 0);
    signal IMF3_9340 : std_logic_vector(7 downto 0);
    signal IMG0_9348 : std_logic_vector(7 downto 0);
    signal IMG1_9356 : std_logic_vector(7 downto 0);
    signal konst_7071_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7081_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7091_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7101_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7111_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7121_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7131_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7141_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7151_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7161_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7171_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7181_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7191_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7201_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7211_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7221_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7231_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7241_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7251_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7261_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7271_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7281_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7291_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7301_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7311_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7321_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7331_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7341_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7351_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7361_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7371_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7381_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7391_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7401_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7411_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7421_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7431_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7441_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7451_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7461_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7471_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7481_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7491_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7501_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7511_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7521_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7531_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7541_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7551_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7561_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7571_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7581_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7591_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7601_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7611_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7621_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7631_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7641_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7651_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7661_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7671_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7681_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7691_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7701_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7711_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7721_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7731_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7741_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7751_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7761_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7771_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7781_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7791_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7801_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7811_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7821_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7831_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7841_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7851_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7861_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7871_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7881_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7891_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7901_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7911_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7921_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7931_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7941_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7951_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7961_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7971_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7981_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7991_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8001_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8011_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8021_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8031_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8041_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8051_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8061_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8071_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8081_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8091_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8101_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8111_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8121_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8131_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8141_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8151_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8161_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8171_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8181_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8191_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8201_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8211_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8221_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8231_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8241_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8251_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8261_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8271_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8281_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8291_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8301_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8311_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8321_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8331_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8341_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8351_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8359_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8367_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8375_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8383_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8391_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8399_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8407_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8415_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8423_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8431_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8439_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8447_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8455_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8463_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8471_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8479_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8487_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8495_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8503_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8511_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8519_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8527_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8535_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8543_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8551_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8559_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8567_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8575_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8583_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8591_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8599_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8607_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8615_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8623_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8631_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8639_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8647_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8655_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8663_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8671_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8679_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8687_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8695_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8703_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8711_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8719_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8727_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8735_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8743_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8751_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8759_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8767_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8775_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8783_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8791_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8799_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8807_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8815_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8823_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8831_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8839_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8847_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8855_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8863_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8871_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8879_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8887_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8895_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8903_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8911_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8919_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8927_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8935_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8943_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8951_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8959_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8967_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8975_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8983_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8991_wire_constant : std_logic_vector(7 downto 0);
    signal konst_8999_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9007_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9015_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9023_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9031_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9039_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9047_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9055_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9063_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9071_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9079_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9087_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9095_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9103_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9111_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9119_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9127_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9135_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9143_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9151_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9159_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9167_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9175_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9183_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9191_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9199_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9207_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9215_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9223_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9231_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9239_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9247_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9255_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9263_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9271_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9279_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9287_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9295_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9303_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9311_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9319_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9327_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9335_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9343_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9351_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9359_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7074_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7076_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7084_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7086_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7094_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7096_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7104_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7106_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7114_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7116_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7124_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7126_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7134_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7136_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7144_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7146_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7154_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7156_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7164_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7166_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7174_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7176_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7184_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7186_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7194_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7196_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7204_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7206_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7214_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7216_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7224_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7226_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7234_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7236_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7244_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7246_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7254_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7256_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7264_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7266_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7274_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7276_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7284_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7286_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7294_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7296_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7304_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7306_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7314_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7316_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7324_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7326_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7334_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7336_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7344_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7346_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7354_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7356_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7364_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7366_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7374_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7376_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7384_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7386_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7394_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7396_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7404_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7406_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7414_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7416_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7424_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7426_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7434_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7436_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7444_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7446_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7454_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7456_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7464_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7466_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7474_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7476_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7484_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7486_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7494_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7496_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7504_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7506_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7514_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7516_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7524_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7526_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7534_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7536_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7544_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7546_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7554_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7556_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7564_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7566_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7574_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7576_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7584_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7586_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7594_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7596_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7604_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7606_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7614_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7616_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7624_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7626_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7634_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7636_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7644_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7646_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7654_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7656_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7664_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7666_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7674_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7676_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7684_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7686_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7694_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7696_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7704_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7706_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7714_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7716_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7724_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7726_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7734_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7736_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7744_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7746_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7754_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7756_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7764_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7766_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7774_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7776_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7784_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7786_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7794_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7796_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7804_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7806_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7814_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7816_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7824_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7826_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7834_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7836_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7844_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7846_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7854_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7856_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7864_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7866_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7874_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7876_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7884_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7886_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7894_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7896_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7904_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7906_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7914_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7916_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7924_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7926_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7934_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7936_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7944_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7946_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7954_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7956_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7964_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7966_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7974_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7976_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7984_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7986_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7994_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_7996_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_8004_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_8006_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_8014_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_8016_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_8024_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_8026_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_8034_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_8036_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_8044_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_8046_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_8054_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_8056_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_8064_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_8066_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_8074_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_8076_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_8084_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_8086_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_8094_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_8096_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_8104_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_8106_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_8114_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_8116_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_8124_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_8126_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_8134_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_8136_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_8144_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_8146_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_8154_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_8156_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_8164_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_8166_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_8174_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_8176_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_8184_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_8186_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_8194_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_8196_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_8204_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_8206_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_8214_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_8216_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_8224_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_8226_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_8234_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_8236_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_8244_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_8246_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_8254_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_8256_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_8264_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_8266_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_8274_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_8276_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_8284_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_8286_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_8294_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_8296_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_8304_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_8306_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_8314_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_8316_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_8324_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_8326_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_8334_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_8336_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_8344_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_8346_wire_constant : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    konst_7071_wire_constant <= "00000000";
    konst_7081_wire_constant <= "00000000";
    konst_7091_wire_constant <= "00000000";
    konst_7101_wire_constant <= "00000000";
    konst_7111_wire_constant <= "00000000";
    konst_7121_wire_constant <= "00000000";
    konst_7131_wire_constant <= "00000000";
    konst_7141_wire_constant <= "00000000";
    konst_7151_wire_constant <= "00000000";
    konst_7161_wire_constant <= "00000000";
    konst_7171_wire_constant <= "00000000";
    konst_7181_wire_constant <= "00000000";
    konst_7191_wire_constant <= "00000000";
    konst_7201_wire_constant <= "00000000";
    konst_7211_wire_constant <= "00000000";
    konst_7221_wire_constant <= "00000000";
    konst_7231_wire_constant <= "00000000";
    konst_7241_wire_constant <= "00000000";
    konst_7251_wire_constant <= "00000000";
    konst_7261_wire_constant <= "00000000";
    konst_7271_wire_constant <= "00000000";
    konst_7281_wire_constant <= "00000000";
    konst_7291_wire_constant <= "00000000";
    konst_7301_wire_constant <= "00000000";
    konst_7311_wire_constant <= "00000000";
    konst_7321_wire_constant <= "00000000";
    konst_7331_wire_constant <= "00000000";
    konst_7341_wire_constant <= "00000000";
    konst_7351_wire_constant <= "00000000";
    konst_7361_wire_constant <= "00000000";
    konst_7371_wire_constant <= "00000000";
    konst_7381_wire_constant <= "00000000";
    konst_7391_wire_constant <= "00000000";
    konst_7401_wire_constant <= "00000000";
    konst_7411_wire_constant <= "00000000";
    konst_7421_wire_constant <= "00000000";
    konst_7431_wire_constant <= "00000000";
    konst_7441_wire_constant <= "00000000";
    konst_7451_wire_constant <= "00000000";
    konst_7461_wire_constant <= "00000000";
    konst_7471_wire_constant <= "00000000";
    konst_7481_wire_constant <= "00000000";
    konst_7491_wire_constant <= "00000000";
    konst_7501_wire_constant <= "00000000";
    konst_7511_wire_constant <= "00000000";
    konst_7521_wire_constant <= "00000000";
    konst_7531_wire_constant <= "00000000";
    konst_7541_wire_constant <= "00000000";
    konst_7551_wire_constant <= "00000000";
    konst_7561_wire_constant <= "00000000";
    konst_7571_wire_constant <= "00000000";
    konst_7581_wire_constant <= "00000000";
    konst_7591_wire_constant <= "00000000";
    konst_7601_wire_constant <= "00000000";
    konst_7611_wire_constant <= "00000000";
    konst_7621_wire_constant <= "00000000";
    konst_7631_wire_constant <= "00000000";
    konst_7641_wire_constant <= "00000000";
    konst_7651_wire_constant <= "00000000";
    konst_7661_wire_constant <= "00000000";
    konst_7671_wire_constant <= "00000000";
    konst_7681_wire_constant <= "00000000";
    konst_7691_wire_constant <= "00000000";
    konst_7701_wire_constant <= "00000000";
    konst_7711_wire_constant <= "00000000";
    konst_7721_wire_constant <= "00000000";
    konst_7731_wire_constant <= "00000000";
    konst_7741_wire_constant <= "00000000";
    konst_7751_wire_constant <= "00000000";
    konst_7761_wire_constant <= "00000000";
    konst_7771_wire_constant <= "00000000";
    konst_7781_wire_constant <= "00000000";
    konst_7791_wire_constant <= "00000000";
    konst_7801_wire_constant <= "00000000";
    konst_7811_wire_constant <= "00000000";
    konst_7821_wire_constant <= "00000000";
    konst_7831_wire_constant <= "00000000";
    konst_7841_wire_constant <= "00000000";
    konst_7851_wire_constant <= "00000000";
    konst_7861_wire_constant <= "00000000";
    konst_7871_wire_constant <= "00000000";
    konst_7881_wire_constant <= "00000000";
    konst_7891_wire_constant <= "00000000";
    konst_7901_wire_constant <= "00000000";
    konst_7911_wire_constant <= "00000000";
    konst_7921_wire_constant <= "00000000";
    konst_7931_wire_constant <= "00000000";
    konst_7941_wire_constant <= "00000000";
    konst_7951_wire_constant <= "00000000";
    konst_7961_wire_constant <= "00000000";
    konst_7971_wire_constant <= "00000000";
    konst_7981_wire_constant <= "00000000";
    konst_7991_wire_constant <= "00000000";
    konst_8001_wire_constant <= "00000000";
    konst_8011_wire_constant <= "00000000";
    konst_8021_wire_constant <= "00000000";
    konst_8031_wire_constant <= "00000000";
    konst_8041_wire_constant <= "00000000";
    konst_8051_wire_constant <= "00000000";
    konst_8061_wire_constant <= "00000000";
    konst_8071_wire_constant <= "00000000";
    konst_8081_wire_constant <= "00000000";
    konst_8091_wire_constant <= "00000000";
    konst_8101_wire_constant <= "00000000";
    konst_8111_wire_constant <= "00000000";
    konst_8121_wire_constant <= "00000000";
    konst_8131_wire_constant <= "00000000";
    konst_8141_wire_constant <= "00000000";
    konst_8151_wire_constant <= "00000000";
    konst_8161_wire_constant <= "00000000";
    konst_8171_wire_constant <= "00000000";
    konst_8181_wire_constant <= "00000000";
    konst_8191_wire_constant <= "00000000";
    konst_8201_wire_constant <= "00000000";
    konst_8211_wire_constant <= "00000000";
    konst_8221_wire_constant <= "00000000";
    konst_8231_wire_constant <= "00000000";
    konst_8241_wire_constant <= "00000000";
    konst_8251_wire_constant <= "00000000";
    konst_8261_wire_constant <= "00000000";
    konst_8271_wire_constant <= "00000000";
    konst_8281_wire_constant <= "00000000";
    konst_8291_wire_constant <= "00000000";
    konst_8301_wire_constant <= "00000000";
    konst_8311_wire_constant <= "00000000";
    konst_8321_wire_constant <= "00000000";
    konst_8331_wire_constant <= "00000000";
    konst_8341_wire_constant <= "00000000";
    konst_8351_wire_constant <= "00000001";
    konst_8359_wire_constant <= "00000001";
    konst_8367_wire_constant <= "00000001";
    konst_8375_wire_constant <= "00000001";
    konst_8383_wire_constant <= "00000001";
    konst_8391_wire_constant <= "00000001";
    konst_8399_wire_constant <= "00000001";
    konst_8407_wire_constant <= "00000001";
    konst_8415_wire_constant <= "00000001";
    konst_8423_wire_constant <= "00000001";
    konst_8431_wire_constant <= "00000001";
    konst_8439_wire_constant <= "00000001";
    konst_8447_wire_constant <= "00000001";
    konst_8455_wire_constant <= "00000001";
    konst_8463_wire_constant <= "00000001";
    konst_8471_wire_constant <= "00000001";
    konst_8479_wire_constant <= "00000001";
    konst_8487_wire_constant <= "00000001";
    konst_8495_wire_constant <= "00000001";
    konst_8503_wire_constant <= "00000001";
    konst_8511_wire_constant <= "00000001";
    konst_8519_wire_constant <= "00000001";
    konst_8527_wire_constant <= "00000001";
    konst_8535_wire_constant <= "00000001";
    konst_8543_wire_constant <= "00000001";
    konst_8551_wire_constant <= "00000001";
    konst_8559_wire_constant <= "00000001";
    konst_8567_wire_constant <= "00000001";
    konst_8575_wire_constant <= "00000001";
    konst_8583_wire_constant <= "00000001";
    konst_8591_wire_constant <= "00000001";
    konst_8599_wire_constant <= "00000001";
    konst_8607_wire_constant <= "00000001";
    konst_8615_wire_constant <= "00000001";
    konst_8623_wire_constant <= "00000001";
    konst_8631_wire_constant <= "00000001";
    konst_8639_wire_constant <= "00000001";
    konst_8647_wire_constant <= "00000001";
    konst_8655_wire_constant <= "00000001";
    konst_8663_wire_constant <= "00000001";
    konst_8671_wire_constant <= "00000001";
    konst_8679_wire_constant <= "00000001";
    konst_8687_wire_constant <= "00000001";
    konst_8695_wire_constant <= "00000001";
    konst_8703_wire_constant <= "00000001";
    konst_8711_wire_constant <= "00000001";
    konst_8719_wire_constant <= "00000001";
    konst_8727_wire_constant <= "00000001";
    konst_8735_wire_constant <= "00000001";
    konst_8743_wire_constant <= "00000001";
    konst_8751_wire_constant <= "00000001";
    konst_8759_wire_constant <= "00000001";
    konst_8767_wire_constant <= "00000001";
    konst_8775_wire_constant <= "00000001";
    konst_8783_wire_constant <= "00000001";
    konst_8791_wire_constant <= "00000001";
    konst_8799_wire_constant <= "00000001";
    konst_8807_wire_constant <= "00000001";
    konst_8815_wire_constant <= "00000001";
    konst_8823_wire_constant <= "00000001";
    konst_8831_wire_constant <= "00000001";
    konst_8839_wire_constant <= "00000001";
    konst_8847_wire_constant <= "00000001";
    konst_8855_wire_constant <= "00000001";
    konst_8863_wire_constant <= "00000010";
    konst_8871_wire_constant <= "00000010";
    konst_8879_wire_constant <= "00000010";
    konst_8887_wire_constant <= "00000010";
    konst_8895_wire_constant <= "00000010";
    konst_8903_wire_constant <= "00000010";
    konst_8911_wire_constant <= "00000010";
    konst_8919_wire_constant <= "00000010";
    konst_8927_wire_constant <= "00000010";
    konst_8935_wire_constant <= "00000010";
    konst_8943_wire_constant <= "00000010";
    konst_8951_wire_constant <= "00000010";
    konst_8959_wire_constant <= "00000010";
    konst_8967_wire_constant <= "00000010";
    konst_8975_wire_constant <= "00000010";
    konst_8983_wire_constant <= "00000010";
    konst_8991_wire_constant <= "00000010";
    konst_8999_wire_constant <= "00000010";
    konst_9007_wire_constant <= "00000010";
    konst_9015_wire_constant <= "00000010";
    konst_9023_wire_constant <= "00000010";
    konst_9031_wire_constant <= "00000010";
    konst_9039_wire_constant <= "00000010";
    konst_9047_wire_constant <= "00000010";
    konst_9055_wire_constant <= "00000010";
    konst_9063_wire_constant <= "00000010";
    konst_9071_wire_constant <= "00000010";
    konst_9079_wire_constant <= "00000010";
    konst_9087_wire_constant <= "00000010";
    konst_9095_wire_constant <= "00000010";
    konst_9103_wire_constant <= "00000010";
    konst_9111_wire_constant <= "00000010";
    konst_9119_wire_constant <= "00000011";
    konst_9127_wire_constant <= "00000011";
    konst_9135_wire_constant <= "00000011";
    konst_9143_wire_constant <= "00000011";
    konst_9151_wire_constant <= "00000011";
    konst_9159_wire_constant <= "00000011";
    konst_9167_wire_constant <= "00000011";
    konst_9175_wire_constant <= "00000011";
    konst_9183_wire_constant <= "00000011";
    konst_9191_wire_constant <= "00000011";
    konst_9199_wire_constant <= "00000011";
    konst_9207_wire_constant <= "00000011";
    konst_9215_wire_constant <= "00000011";
    konst_9223_wire_constant <= "00000011";
    konst_9231_wire_constant <= "00000011";
    konst_9239_wire_constant <= "00000011";
    konst_9247_wire_constant <= "00000100";
    konst_9255_wire_constant <= "00000100";
    konst_9263_wire_constant <= "00000100";
    konst_9271_wire_constant <= "00000100";
    konst_9279_wire_constant <= "00000100";
    konst_9287_wire_constant <= "00000100";
    konst_9295_wire_constant <= "00000100";
    konst_9303_wire_constant <= "00000100";
    konst_9311_wire_constant <= "00000101";
    konst_9319_wire_constant <= "00000101";
    konst_9327_wire_constant <= "00000101";
    konst_9335_wire_constant <= "00000101";
    konst_9343_wire_constant <= "00000110";
    konst_9351_wire_constant <= "00000110";
    konst_9359_wire_constant <= "00000111";
    type_cast_7074_wire_constant <= "00001001";
    type_cast_7076_wire_constant <= "01010010";
    type_cast_7084_wire_constant <= "11010101";
    type_cast_7086_wire_constant <= "01101010";
    type_cast_7094_wire_constant <= "00110110";
    type_cast_7096_wire_constant <= "00110000";
    type_cast_7104_wire_constant <= "00111000";
    type_cast_7106_wire_constant <= "10100101";
    type_cast_7114_wire_constant <= "01000000";
    type_cast_7116_wire_constant <= "10111111";
    type_cast_7124_wire_constant <= "10011110";
    type_cast_7126_wire_constant <= "10100011";
    type_cast_7134_wire_constant <= "11110011";
    type_cast_7136_wire_constant <= "10000001";
    type_cast_7144_wire_constant <= "11111011";
    type_cast_7146_wire_constant <= "11010111";
    type_cast_7154_wire_constant <= "11100011";
    type_cast_7156_wire_constant <= "01111100";
    type_cast_7164_wire_constant <= "10000010";
    type_cast_7166_wire_constant <= "00111001";
    type_cast_7174_wire_constant <= "00101111";
    type_cast_7176_wire_constant <= "10011011";
    type_cast_7184_wire_constant <= "10000111";
    type_cast_7186_wire_constant <= "11111111";
    type_cast_7194_wire_constant <= "10001110";
    type_cast_7196_wire_constant <= "00110100";
    type_cast_7204_wire_constant <= "01000100";
    type_cast_7206_wire_constant <= "01000011";
    type_cast_7214_wire_constant <= "11011110";
    type_cast_7216_wire_constant <= "11000100";
    type_cast_7224_wire_constant <= "11001011";
    type_cast_7226_wire_constant <= "11101001";
    type_cast_7234_wire_constant <= "01111011";
    type_cast_7236_wire_constant <= "01010100";
    type_cast_7244_wire_constant <= "00110010";
    type_cast_7246_wire_constant <= "10010100";
    type_cast_7254_wire_constant <= "11000010";
    type_cast_7256_wire_constant <= "10100110";
    type_cast_7264_wire_constant <= "00111101";
    type_cast_7266_wire_constant <= "00100011";
    type_cast_7274_wire_constant <= "01001100";
    type_cast_7276_wire_constant <= "11101110";
    type_cast_7284_wire_constant <= "00001011";
    type_cast_7286_wire_constant <= "10010101";
    type_cast_7294_wire_constant <= "11111010";
    type_cast_7296_wire_constant <= "01000010";
    type_cast_7304_wire_constant <= "01001110";
    type_cast_7306_wire_constant <= "11000011";
    type_cast_7314_wire_constant <= "00101110";
    type_cast_7316_wire_constant <= "00001000";
    type_cast_7324_wire_constant <= "01100110";
    type_cast_7326_wire_constant <= "10100001";
    type_cast_7334_wire_constant <= "11011001";
    type_cast_7336_wire_constant <= "00101000";
    type_cast_7344_wire_constant <= "10110010";
    type_cast_7346_wire_constant <= "00100100";
    type_cast_7354_wire_constant <= "01011011";
    type_cast_7356_wire_constant <= "01110110";
    type_cast_7364_wire_constant <= "01001001";
    type_cast_7366_wire_constant <= "10100010";
    type_cast_7374_wire_constant <= "10001011";
    type_cast_7376_wire_constant <= "01101101";
    type_cast_7384_wire_constant <= "00100101";
    type_cast_7386_wire_constant <= "11010001";
    type_cast_7394_wire_constant <= "11111000";
    type_cast_7396_wire_constant <= "01110010";
    type_cast_7404_wire_constant <= "01100100";
    type_cast_7406_wire_constant <= "11110110";
    type_cast_7414_wire_constant <= "01101000";
    type_cast_7416_wire_constant <= "10000110";
    type_cast_7424_wire_constant <= "00010110";
    type_cast_7426_wire_constant <= "10011000";
    type_cast_7434_wire_constant <= "10100100";
    type_cast_7436_wire_constant <= "11010100";
    type_cast_7444_wire_constant <= "11001100";
    type_cast_7446_wire_constant <= "01011100";
    type_cast_7454_wire_constant <= "01100101";
    type_cast_7456_wire_constant <= "01011101";
    type_cast_7464_wire_constant <= "10010010";
    type_cast_7466_wire_constant <= "10110110";
    type_cast_7474_wire_constant <= "01110000";
    type_cast_7476_wire_constant <= "01101100";
    type_cast_7484_wire_constant <= "01010000";
    type_cast_7486_wire_constant <= "01001000";
    type_cast_7494_wire_constant <= "11101101";
    type_cast_7496_wire_constant <= "11111101";
    type_cast_7504_wire_constant <= "11011010";
    type_cast_7506_wire_constant <= "10111001";
    type_cast_7514_wire_constant <= "00010101";
    type_cast_7516_wire_constant <= "01011110";
    type_cast_7524_wire_constant <= "01010111";
    type_cast_7526_wire_constant <= "01000110";
    type_cast_7534_wire_constant <= "10001101";
    type_cast_7536_wire_constant <= "10100111";
    type_cast_7544_wire_constant <= "10000100";
    type_cast_7546_wire_constant <= "10011101";
    type_cast_7554_wire_constant <= "11011000";
    type_cast_7556_wire_constant <= "10010000";
    type_cast_7564_wire_constant <= "00000000";
    type_cast_7566_wire_constant <= "10101011";
    type_cast_7574_wire_constant <= "10111100";
    type_cast_7576_wire_constant <= "10001100";
    type_cast_7584_wire_constant <= "00001010";
    type_cast_7586_wire_constant <= "11010011";
    type_cast_7594_wire_constant <= "11100100";
    type_cast_7596_wire_constant <= "11110111";
    type_cast_7604_wire_constant <= "00000101";
    type_cast_7606_wire_constant <= "01011000";
    type_cast_7614_wire_constant <= "10110011";
    type_cast_7616_wire_constant <= "10111000";
    type_cast_7624_wire_constant <= "00000110";
    type_cast_7626_wire_constant <= "01000101";
    type_cast_7634_wire_constant <= "00101100";
    type_cast_7636_wire_constant <= "11010000";
    type_cast_7644_wire_constant <= "10001111";
    type_cast_7646_wire_constant <= "00011110";
    type_cast_7654_wire_constant <= "00111111";
    type_cast_7656_wire_constant <= "11001010";
    type_cast_7664_wire_constant <= "00000010";
    type_cast_7666_wire_constant <= "00001111";
    type_cast_7674_wire_constant <= "10101111";
    type_cast_7676_wire_constant <= "11000001";
    type_cast_7684_wire_constant <= "00000011";
    type_cast_7686_wire_constant <= "10111101";
    type_cast_7694_wire_constant <= "00010011";
    type_cast_7696_wire_constant <= "00000001";
    type_cast_7704_wire_constant <= "01101011";
    type_cast_7706_wire_constant <= "10001010";
    type_cast_7714_wire_constant <= "10010001";
    type_cast_7716_wire_constant <= "00111010";
    type_cast_7724_wire_constant <= "01000001";
    type_cast_7726_wire_constant <= "00010001";
    type_cast_7734_wire_constant <= "01100111";
    type_cast_7736_wire_constant <= "01001111";
    type_cast_7744_wire_constant <= "11101010";
    type_cast_7746_wire_constant <= "11011100";
    type_cast_7754_wire_constant <= "11110010";
    type_cast_7756_wire_constant <= "10010111";
    type_cast_7764_wire_constant <= "11001110";
    type_cast_7766_wire_constant <= "11001111";
    type_cast_7774_wire_constant <= "10110100";
    type_cast_7776_wire_constant <= "11110000";
    type_cast_7784_wire_constant <= "01110011";
    type_cast_7786_wire_constant <= "11100110";
    type_cast_7794_wire_constant <= "10101100";
    type_cast_7796_wire_constant <= "10010110";
    type_cast_7804_wire_constant <= "00100010";
    type_cast_7806_wire_constant <= "01110100";
    type_cast_7814_wire_constant <= "10101101";
    type_cast_7816_wire_constant <= "11100111";
    type_cast_7824_wire_constant <= "10000101";
    type_cast_7826_wire_constant <= "00110101";
    type_cast_7834_wire_constant <= "11111001";
    type_cast_7836_wire_constant <= "11100010";
    type_cast_7844_wire_constant <= "11101000";
    type_cast_7846_wire_constant <= "00110111";
    type_cast_7854_wire_constant <= "01110101";
    type_cast_7856_wire_constant <= "00011100";
    type_cast_7864_wire_constant <= "01101110";
    type_cast_7866_wire_constant <= "11011111";
    type_cast_7874_wire_constant <= "11110001";
    type_cast_7876_wire_constant <= "01000111";
    type_cast_7884_wire_constant <= "01110001";
    type_cast_7886_wire_constant <= "00011010";
    type_cast_7894_wire_constant <= "00101001";
    type_cast_7896_wire_constant <= "00011101";
    type_cast_7904_wire_constant <= "10001001";
    type_cast_7906_wire_constant <= "11000101";
    type_cast_7914_wire_constant <= "10110111";
    type_cast_7916_wire_constant <= "01101111";
    type_cast_7924_wire_constant <= "00001110";
    type_cast_7926_wire_constant <= "01100010";
    type_cast_7934_wire_constant <= "00011000";
    type_cast_7936_wire_constant <= "10101010";
    type_cast_7944_wire_constant <= "00011011";
    type_cast_7946_wire_constant <= "10111110";
    type_cast_7954_wire_constant <= "01010110";
    type_cast_7956_wire_constant <= "11111100";
    type_cast_7964_wire_constant <= "01001011";
    type_cast_7966_wire_constant <= "00111110";
    type_cast_7974_wire_constant <= "11010010";
    type_cast_7976_wire_constant <= "11000110";
    type_cast_7984_wire_constant <= "00100000";
    type_cast_7986_wire_constant <= "01111001";
    type_cast_7994_wire_constant <= "11011011";
    type_cast_7996_wire_constant <= "10011010";
    type_cast_8004_wire_constant <= "11111110";
    type_cast_8006_wire_constant <= "11000000";
    type_cast_8014_wire_constant <= "11001101";
    type_cast_8016_wire_constant <= "01111000";
    type_cast_8024_wire_constant <= "11110100";
    type_cast_8026_wire_constant <= "01011010";
    type_cast_8034_wire_constant <= "11011101";
    type_cast_8036_wire_constant <= "00011111";
    type_cast_8044_wire_constant <= "00110011";
    type_cast_8046_wire_constant <= "10101000";
    type_cast_8054_wire_constant <= "00000111";
    type_cast_8056_wire_constant <= "10001000";
    type_cast_8064_wire_constant <= "00110001";
    type_cast_8066_wire_constant <= "11000111";
    type_cast_8074_wire_constant <= "00010010";
    type_cast_8076_wire_constant <= "10110001";
    type_cast_8084_wire_constant <= "01011001";
    type_cast_8086_wire_constant <= "00010000";
    type_cast_8094_wire_constant <= "10000000";
    type_cast_8096_wire_constant <= "00100111";
    type_cast_8104_wire_constant <= "01011111";
    type_cast_8106_wire_constant <= "11101100";
    type_cast_8114_wire_constant <= "01010001";
    type_cast_8116_wire_constant <= "01100000";
    type_cast_8124_wire_constant <= "10101001";
    type_cast_8126_wire_constant <= "01111111";
    type_cast_8134_wire_constant <= "10110101";
    type_cast_8136_wire_constant <= "00011001";
    type_cast_8144_wire_constant <= "00001101";
    type_cast_8146_wire_constant <= "01001010";
    type_cast_8154_wire_constant <= "11100101";
    type_cast_8156_wire_constant <= "00101101";
    type_cast_8164_wire_constant <= "10011111";
    type_cast_8166_wire_constant <= "01111010";
    type_cast_8174_wire_constant <= "11001001";
    type_cast_8176_wire_constant <= "10010011";
    type_cast_8184_wire_constant <= "11101111";
    type_cast_8186_wire_constant <= "10011100";
    type_cast_8194_wire_constant <= "11100000";
    type_cast_8196_wire_constant <= "10100000";
    type_cast_8204_wire_constant <= "01001101";
    type_cast_8206_wire_constant <= "00111011";
    type_cast_8214_wire_constant <= "00101010";
    type_cast_8216_wire_constant <= "10101110";
    type_cast_8224_wire_constant <= "10110000";
    type_cast_8226_wire_constant <= "11110101";
    type_cast_8234_wire_constant <= "11101011";
    type_cast_8236_wire_constant <= "11001000";
    type_cast_8244_wire_constant <= "00111100";
    type_cast_8246_wire_constant <= "10111011";
    type_cast_8254_wire_constant <= "01010011";
    type_cast_8256_wire_constant <= "10000011";
    type_cast_8264_wire_constant <= "01100001";
    type_cast_8266_wire_constant <= "10011001";
    type_cast_8274_wire_constant <= "00101011";
    type_cast_8276_wire_constant <= "00010111";
    type_cast_8284_wire_constant <= "01111110";
    type_cast_8286_wire_constant <= "00000100";
    type_cast_8294_wire_constant <= "01110111";
    type_cast_8296_wire_constant <= "10111010";
    type_cast_8304_wire_constant <= "00100110";
    type_cast_8306_wire_constant <= "11010110";
    type_cast_8314_wire_constant <= "01101001";
    type_cast_8316_wire_constant <= "11100001";
    type_cast_8324_wire_constant <= "01100011";
    type_cast_8326_wire_constant <= "00010100";
    type_cast_8334_wire_constant <= "00100001";
    type_cast_8336_wire_constant <= "01010101";
    type_cast_8344_wire_constant <= "01111101";
    type_cast_8346_wire_constant <= "00001100";
    -- flow-through select operator MUX_7077_inst
    IMA0_7078 <= type_cast_7074_wire_constant when (BITSEL_u8_u1_7072_wire(0) /=  '0') else type_cast_7076_wire_constant;
    -- flow-through select operator MUX_7087_inst
    IMA1_7088 <= type_cast_7084_wire_constant when (BITSEL_u8_u1_7082_wire(0) /=  '0') else type_cast_7086_wire_constant;
    -- flow-through select operator MUX_7097_inst
    IMA2_7098 <= type_cast_7094_wire_constant when (BITSEL_u8_u1_7092_wire(0) /=  '0') else type_cast_7096_wire_constant;
    -- flow-through select operator MUX_7107_inst
    IMA3_7108 <= type_cast_7104_wire_constant when (BITSEL_u8_u1_7102_wire(0) /=  '0') else type_cast_7106_wire_constant;
    -- flow-through select operator MUX_7117_inst
    IMA4_7118 <= type_cast_7114_wire_constant when (BITSEL_u8_u1_7112_wire(0) /=  '0') else type_cast_7116_wire_constant;
    -- flow-through select operator MUX_7127_inst
    IMA5_7128 <= type_cast_7124_wire_constant when (BITSEL_u8_u1_7122_wire(0) /=  '0') else type_cast_7126_wire_constant;
    -- flow-through select operator MUX_7137_inst
    IMA6_7138 <= type_cast_7134_wire_constant when (BITSEL_u8_u1_7132_wire(0) /=  '0') else type_cast_7136_wire_constant;
    -- flow-through select operator MUX_7147_inst
    IMA7_7148 <= type_cast_7144_wire_constant when (BITSEL_u8_u1_7142_wire(0) /=  '0') else type_cast_7146_wire_constant;
    -- flow-through select operator MUX_7157_inst
    IMA8_7158 <= type_cast_7154_wire_constant when (BITSEL_u8_u1_7152_wire(0) /=  '0') else type_cast_7156_wire_constant;
    -- flow-through select operator MUX_7167_inst
    IMA9_7168 <= type_cast_7164_wire_constant when (BITSEL_u8_u1_7162_wire(0) /=  '0') else type_cast_7166_wire_constant;
    -- flow-through select operator MUX_7177_inst
    IMA10_7178 <= type_cast_7174_wire_constant when (BITSEL_u8_u1_7172_wire(0) /=  '0') else type_cast_7176_wire_constant;
    -- flow-through select operator MUX_7187_inst
    IMA11_7188 <= type_cast_7184_wire_constant when (BITSEL_u8_u1_7182_wire(0) /=  '0') else type_cast_7186_wire_constant;
    -- flow-through select operator MUX_7197_inst
    IMA12_7198 <= type_cast_7194_wire_constant when (BITSEL_u8_u1_7192_wire(0) /=  '0') else type_cast_7196_wire_constant;
    -- flow-through select operator MUX_7207_inst
    IMA13_7208 <= type_cast_7204_wire_constant when (BITSEL_u8_u1_7202_wire(0) /=  '0') else type_cast_7206_wire_constant;
    -- flow-through select operator MUX_7217_inst
    IMA14_7218 <= type_cast_7214_wire_constant when (BITSEL_u8_u1_7212_wire(0) /=  '0') else type_cast_7216_wire_constant;
    -- flow-through select operator MUX_7227_inst
    IMA15_7228 <= type_cast_7224_wire_constant when (BITSEL_u8_u1_7222_wire(0) /=  '0') else type_cast_7226_wire_constant;
    -- flow-through select operator MUX_7237_inst
    IMA16_7238 <= type_cast_7234_wire_constant when (BITSEL_u8_u1_7232_wire(0) /=  '0') else type_cast_7236_wire_constant;
    -- flow-through select operator MUX_7247_inst
    IMA17_7248 <= type_cast_7244_wire_constant when (BITSEL_u8_u1_7242_wire(0) /=  '0') else type_cast_7246_wire_constant;
    -- flow-through select operator MUX_7257_inst
    IMA18_7258 <= type_cast_7254_wire_constant when (BITSEL_u8_u1_7252_wire(0) /=  '0') else type_cast_7256_wire_constant;
    -- flow-through select operator MUX_7267_inst
    IMA19_7268 <= type_cast_7264_wire_constant when (BITSEL_u8_u1_7262_wire(0) /=  '0') else type_cast_7266_wire_constant;
    -- flow-through select operator MUX_7277_inst
    IMA20_7278 <= type_cast_7274_wire_constant when (BITSEL_u8_u1_7272_wire(0) /=  '0') else type_cast_7276_wire_constant;
    -- flow-through select operator MUX_7287_inst
    IMA21_7288 <= type_cast_7284_wire_constant when (BITSEL_u8_u1_7282_wire(0) /=  '0') else type_cast_7286_wire_constant;
    -- flow-through select operator MUX_7297_inst
    IMA22_7298 <= type_cast_7294_wire_constant when (BITSEL_u8_u1_7292_wire(0) /=  '0') else type_cast_7296_wire_constant;
    -- flow-through select operator MUX_7307_inst
    IMA23_7308 <= type_cast_7304_wire_constant when (BITSEL_u8_u1_7302_wire(0) /=  '0') else type_cast_7306_wire_constant;
    -- flow-through select operator MUX_7317_inst
    IMA24_7318 <= type_cast_7314_wire_constant when (BITSEL_u8_u1_7312_wire(0) /=  '0') else type_cast_7316_wire_constant;
    -- flow-through select operator MUX_7327_inst
    IMA25_7328 <= type_cast_7324_wire_constant when (BITSEL_u8_u1_7322_wire(0) /=  '0') else type_cast_7326_wire_constant;
    -- flow-through select operator MUX_7337_inst
    IMA26_7338 <= type_cast_7334_wire_constant when (BITSEL_u8_u1_7332_wire(0) /=  '0') else type_cast_7336_wire_constant;
    -- flow-through select operator MUX_7347_inst
    IMA27_7348 <= type_cast_7344_wire_constant when (BITSEL_u8_u1_7342_wire(0) /=  '0') else type_cast_7346_wire_constant;
    -- flow-through select operator MUX_7357_inst
    IMA28_7358 <= type_cast_7354_wire_constant when (BITSEL_u8_u1_7352_wire(0) /=  '0') else type_cast_7356_wire_constant;
    -- flow-through select operator MUX_7367_inst
    IMA29_7368 <= type_cast_7364_wire_constant when (BITSEL_u8_u1_7362_wire(0) /=  '0') else type_cast_7366_wire_constant;
    -- flow-through select operator MUX_7377_inst
    IMA30_7378 <= type_cast_7374_wire_constant when (BITSEL_u8_u1_7372_wire(0) /=  '0') else type_cast_7376_wire_constant;
    -- flow-through select operator MUX_7387_inst
    IMA31_7388 <= type_cast_7384_wire_constant when (BITSEL_u8_u1_7382_wire(0) /=  '0') else type_cast_7386_wire_constant;
    -- flow-through select operator MUX_7397_inst
    IMA32_7398 <= type_cast_7394_wire_constant when (BITSEL_u8_u1_7392_wire(0) /=  '0') else type_cast_7396_wire_constant;
    -- flow-through select operator MUX_7407_inst
    IMA33_7408 <= type_cast_7404_wire_constant when (BITSEL_u8_u1_7402_wire(0) /=  '0') else type_cast_7406_wire_constant;
    -- flow-through select operator MUX_7417_inst
    IMA34_7418 <= type_cast_7414_wire_constant when (BITSEL_u8_u1_7412_wire(0) /=  '0') else type_cast_7416_wire_constant;
    -- flow-through select operator MUX_7427_inst
    IMA35_7428 <= type_cast_7424_wire_constant when (BITSEL_u8_u1_7422_wire(0) /=  '0') else type_cast_7426_wire_constant;
    -- flow-through select operator MUX_7437_inst
    IMA36_7438 <= type_cast_7434_wire_constant when (BITSEL_u8_u1_7432_wire(0) /=  '0') else type_cast_7436_wire_constant;
    -- flow-through select operator MUX_7447_inst
    IMA37_7448 <= type_cast_7444_wire_constant when (BITSEL_u8_u1_7442_wire(0) /=  '0') else type_cast_7446_wire_constant;
    -- flow-through select operator MUX_7457_inst
    IMA38_7458 <= type_cast_7454_wire_constant when (BITSEL_u8_u1_7452_wire(0) /=  '0') else type_cast_7456_wire_constant;
    -- flow-through select operator MUX_7467_inst
    IMA39_7468 <= type_cast_7464_wire_constant when (BITSEL_u8_u1_7462_wire(0) /=  '0') else type_cast_7466_wire_constant;
    -- flow-through select operator MUX_7477_inst
    IMA40_7478 <= type_cast_7474_wire_constant when (BITSEL_u8_u1_7472_wire(0) /=  '0') else type_cast_7476_wire_constant;
    -- flow-through select operator MUX_7487_inst
    IMA41_7488 <= type_cast_7484_wire_constant when (BITSEL_u8_u1_7482_wire(0) /=  '0') else type_cast_7486_wire_constant;
    -- flow-through select operator MUX_7497_inst
    IMA42_7498 <= type_cast_7494_wire_constant when (BITSEL_u8_u1_7492_wire(0) /=  '0') else type_cast_7496_wire_constant;
    -- flow-through select operator MUX_7507_inst
    IMA43_7508 <= type_cast_7504_wire_constant when (BITSEL_u8_u1_7502_wire(0) /=  '0') else type_cast_7506_wire_constant;
    -- flow-through select operator MUX_7517_inst
    IMA44_7518 <= type_cast_7514_wire_constant when (BITSEL_u8_u1_7512_wire(0) /=  '0') else type_cast_7516_wire_constant;
    -- flow-through select operator MUX_7527_inst
    IMA45_7528 <= type_cast_7524_wire_constant when (BITSEL_u8_u1_7522_wire(0) /=  '0') else type_cast_7526_wire_constant;
    -- flow-through select operator MUX_7537_inst
    IMA46_7538 <= type_cast_7534_wire_constant when (BITSEL_u8_u1_7532_wire(0) /=  '0') else type_cast_7536_wire_constant;
    -- flow-through select operator MUX_7547_inst
    IMA47_7548 <= type_cast_7544_wire_constant when (BITSEL_u8_u1_7542_wire(0) /=  '0') else type_cast_7546_wire_constant;
    -- flow-through select operator MUX_7557_inst
    IMA48_7558 <= type_cast_7554_wire_constant when (BITSEL_u8_u1_7552_wire(0) /=  '0') else type_cast_7556_wire_constant;
    -- flow-through select operator MUX_7567_inst
    IMA49_7568 <= type_cast_7564_wire_constant when (BITSEL_u8_u1_7562_wire(0) /=  '0') else type_cast_7566_wire_constant;
    -- flow-through select operator MUX_7577_inst
    IMA50_7578 <= type_cast_7574_wire_constant when (BITSEL_u8_u1_7572_wire(0) /=  '0') else type_cast_7576_wire_constant;
    -- flow-through select operator MUX_7587_inst
    IMA51_7588 <= type_cast_7584_wire_constant when (BITSEL_u8_u1_7582_wire(0) /=  '0') else type_cast_7586_wire_constant;
    -- flow-through select operator MUX_7597_inst
    IMA52_7598 <= type_cast_7594_wire_constant when (BITSEL_u8_u1_7592_wire(0) /=  '0') else type_cast_7596_wire_constant;
    -- flow-through select operator MUX_7607_inst
    IMA53_7608 <= type_cast_7604_wire_constant when (BITSEL_u8_u1_7602_wire(0) /=  '0') else type_cast_7606_wire_constant;
    -- flow-through select operator MUX_7617_inst
    IMA54_7618 <= type_cast_7614_wire_constant when (BITSEL_u8_u1_7612_wire(0) /=  '0') else type_cast_7616_wire_constant;
    -- flow-through select operator MUX_7627_inst
    IMA55_7628 <= type_cast_7624_wire_constant when (BITSEL_u8_u1_7622_wire(0) /=  '0') else type_cast_7626_wire_constant;
    -- flow-through select operator MUX_7637_inst
    IMA56_7638 <= type_cast_7634_wire_constant when (BITSEL_u8_u1_7632_wire(0) /=  '0') else type_cast_7636_wire_constant;
    -- flow-through select operator MUX_7647_inst
    IMA57_7648 <= type_cast_7644_wire_constant when (BITSEL_u8_u1_7642_wire(0) /=  '0') else type_cast_7646_wire_constant;
    -- flow-through select operator MUX_7657_inst
    IMA58_7658 <= type_cast_7654_wire_constant when (BITSEL_u8_u1_7652_wire(0) /=  '0') else type_cast_7656_wire_constant;
    -- flow-through select operator MUX_7667_inst
    IMA59_7668 <= type_cast_7664_wire_constant when (BITSEL_u8_u1_7662_wire(0) /=  '0') else type_cast_7666_wire_constant;
    -- flow-through select operator MUX_7677_inst
    IMA60_7678 <= type_cast_7674_wire_constant when (BITSEL_u8_u1_7672_wire(0) /=  '0') else type_cast_7676_wire_constant;
    -- flow-through select operator MUX_7687_inst
    IMA61_7688 <= type_cast_7684_wire_constant when (BITSEL_u8_u1_7682_wire(0) /=  '0') else type_cast_7686_wire_constant;
    -- flow-through select operator MUX_7697_inst
    IMA62_7698 <= type_cast_7694_wire_constant when (BITSEL_u8_u1_7692_wire(0) /=  '0') else type_cast_7696_wire_constant;
    -- flow-through select operator MUX_7707_inst
    IMA63_7708 <= type_cast_7704_wire_constant when (BITSEL_u8_u1_7702_wire(0) /=  '0') else type_cast_7706_wire_constant;
    -- flow-through select operator MUX_7717_inst
    IMA64_7718 <= type_cast_7714_wire_constant when (BITSEL_u8_u1_7712_wire(0) /=  '0') else type_cast_7716_wire_constant;
    -- flow-through select operator MUX_7727_inst
    IMA65_7728 <= type_cast_7724_wire_constant when (BITSEL_u8_u1_7722_wire(0) /=  '0') else type_cast_7726_wire_constant;
    -- flow-through select operator MUX_7737_inst
    IMA66_7738 <= type_cast_7734_wire_constant when (BITSEL_u8_u1_7732_wire(0) /=  '0') else type_cast_7736_wire_constant;
    -- flow-through select operator MUX_7747_inst
    IMA67_7748 <= type_cast_7744_wire_constant when (BITSEL_u8_u1_7742_wire(0) /=  '0') else type_cast_7746_wire_constant;
    -- flow-through select operator MUX_7757_inst
    IMA68_7758 <= type_cast_7754_wire_constant when (BITSEL_u8_u1_7752_wire(0) /=  '0') else type_cast_7756_wire_constant;
    -- flow-through select operator MUX_7767_inst
    IMA69_7768 <= type_cast_7764_wire_constant when (BITSEL_u8_u1_7762_wire(0) /=  '0') else type_cast_7766_wire_constant;
    -- flow-through select operator MUX_7777_inst
    IMA70_7778 <= type_cast_7774_wire_constant when (BITSEL_u8_u1_7772_wire(0) /=  '0') else type_cast_7776_wire_constant;
    -- flow-through select operator MUX_7787_inst
    IMA71_7788 <= type_cast_7784_wire_constant when (BITSEL_u8_u1_7782_wire(0) /=  '0') else type_cast_7786_wire_constant;
    -- flow-through select operator MUX_7797_inst
    IMA72_7798 <= type_cast_7794_wire_constant when (BITSEL_u8_u1_7792_wire(0) /=  '0') else type_cast_7796_wire_constant;
    -- flow-through select operator MUX_7807_inst
    IMA73_7808 <= type_cast_7804_wire_constant when (BITSEL_u8_u1_7802_wire(0) /=  '0') else type_cast_7806_wire_constant;
    -- flow-through select operator MUX_7817_inst
    IMA74_7818 <= type_cast_7814_wire_constant when (BITSEL_u8_u1_7812_wire(0) /=  '0') else type_cast_7816_wire_constant;
    -- flow-through select operator MUX_7827_inst
    IMA75_7828 <= type_cast_7824_wire_constant when (BITSEL_u8_u1_7822_wire(0) /=  '0') else type_cast_7826_wire_constant;
    -- flow-through select operator MUX_7837_inst
    IMA76_7838 <= type_cast_7834_wire_constant when (BITSEL_u8_u1_7832_wire(0) /=  '0') else type_cast_7836_wire_constant;
    -- flow-through select operator MUX_7847_inst
    IMA77_7848 <= type_cast_7844_wire_constant when (BITSEL_u8_u1_7842_wire(0) /=  '0') else type_cast_7846_wire_constant;
    -- flow-through select operator MUX_7857_inst
    IMA78_7858 <= type_cast_7854_wire_constant when (BITSEL_u8_u1_7852_wire(0) /=  '0') else type_cast_7856_wire_constant;
    -- flow-through select operator MUX_7867_inst
    IMA79_7868 <= type_cast_7864_wire_constant when (BITSEL_u8_u1_7862_wire(0) /=  '0') else type_cast_7866_wire_constant;
    -- flow-through select operator MUX_7877_inst
    IMA80_7878 <= type_cast_7874_wire_constant when (BITSEL_u8_u1_7872_wire(0) /=  '0') else type_cast_7876_wire_constant;
    -- flow-through select operator MUX_7887_inst
    IMA81_7888 <= type_cast_7884_wire_constant when (BITSEL_u8_u1_7882_wire(0) /=  '0') else type_cast_7886_wire_constant;
    -- flow-through select operator MUX_7897_inst
    IMA82_7898 <= type_cast_7894_wire_constant when (BITSEL_u8_u1_7892_wire(0) /=  '0') else type_cast_7896_wire_constant;
    -- flow-through select operator MUX_7907_inst
    IMA83_7908 <= type_cast_7904_wire_constant when (BITSEL_u8_u1_7902_wire(0) /=  '0') else type_cast_7906_wire_constant;
    -- flow-through select operator MUX_7917_inst
    IMA84_7918 <= type_cast_7914_wire_constant when (BITSEL_u8_u1_7912_wire(0) /=  '0') else type_cast_7916_wire_constant;
    -- flow-through select operator MUX_7927_inst
    IMA85_7928 <= type_cast_7924_wire_constant when (BITSEL_u8_u1_7922_wire(0) /=  '0') else type_cast_7926_wire_constant;
    -- flow-through select operator MUX_7937_inst
    IMA86_7938 <= type_cast_7934_wire_constant when (BITSEL_u8_u1_7932_wire(0) /=  '0') else type_cast_7936_wire_constant;
    -- flow-through select operator MUX_7947_inst
    IMA87_7948 <= type_cast_7944_wire_constant when (BITSEL_u8_u1_7942_wire(0) /=  '0') else type_cast_7946_wire_constant;
    -- flow-through select operator MUX_7957_inst
    IMA88_7958 <= type_cast_7954_wire_constant when (BITSEL_u8_u1_7952_wire(0) /=  '0') else type_cast_7956_wire_constant;
    -- flow-through select operator MUX_7967_inst
    IMA89_7968 <= type_cast_7964_wire_constant when (BITSEL_u8_u1_7962_wire(0) /=  '0') else type_cast_7966_wire_constant;
    -- flow-through select operator MUX_7977_inst
    IMA90_7978 <= type_cast_7974_wire_constant when (BITSEL_u8_u1_7972_wire(0) /=  '0') else type_cast_7976_wire_constant;
    -- flow-through select operator MUX_7987_inst
    IMA91_7988 <= type_cast_7984_wire_constant when (BITSEL_u8_u1_7982_wire(0) /=  '0') else type_cast_7986_wire_constant;
    -- flow-through select operator MUX_7997_inst
    IMA92_7998 <= type_cast_7994_wire_constant when (BITSEL_u8_u1_7992_wire(0) /=  '0') else type_cast_7996_wire_constant;
    -- flow-through select operator MUX_8007_inst
    IMA93_8008 <= type_cast_8004_wire_constant when (BITSEL_u8_u1_8002_wire(0) /=  '0') else type_cast_8006_wire_constant;
    -- flow-through select operator MUX_8017_inst
    IMA94_8018 <= type_cast_8014_wire_constant when (BITSEL_u8_u1_8012_wire(0) /=  '0') else type_cast_8016_wire_constant;
    -- flow-through select operator MUX_8027_inst
    IMA95_8028 <= type_cast_8024_wire_constant when (BITSEL_u8_u1_8022_wire(0) /=  '0') else type_cast_8026_wire_constant;
    -- flow-through select operator MUX_8037_inst
    IMA96_8038 <= type_cast_8034_wire_constant when (BITSEL_u8_u1_8032_wire(0) /=  '0') else type_cast_8036_wire_constant;
    -- flow-through select operator MUX_8047_inst
    IMA97_8048 <= type_cast_8044_wire_constant when (BITSEL_u8_u1_8042_wire(0) /=  '0') else type_cast_8046_wire_constant;
    -- flow-through select operator MUX_8057_inst
    IMA98_8058 <= type_cast_8054_wire_constant when (BITSEL_u8_u1_8052_wire(0) /=  '0') else type_cast_8056_wire_constant;
    -- flow-through select operator MUX_8067_inst
    IMA99_8068 <= type_cast_8064_wire_constant when (BITSEL_u8_u1_8062_wire(0) /=  '0') else type_cast_8066_wire_constant;
    -- flow-through select operator MUX_8077_inst
    IMA100_8078 <= type_cast_8074_wire_constant when (BITSEL_u8_u1_8072_wire(0) /=  '0') else type_cast_8076_wire_constant;
    -- flow-through select operator MUX_8087_inst
    IMA101_8088 <= type_cast_8084_wire_constant when (BITSEL_u8_u1_8082_wire(0) /=  '0') else type_cast_8086_wire_constant;
    -- flow-through select operator MUX_8097_inst
    IMA102_8098 <= type_cast_8094_wire_constant when (BITSEL_u8_u1_8092_wire(0) /=  '0') else type_cast_8096_wire_constant;
    -- flow-through select operator MUX_8107_inst
    IMA103_8108 <= type_cast_8104_wire_constant when (BITSEL_u8_u1_8102_wire(0) /=  '0') else type_cast_8106_wire_constant;
    -- flow-through select operator MUX_8117_inst
    IMA104_8118 <= type_cast_8114_wire_constant when (BITSEL_u8_u1_8112_wire(0) /=  '0') else type_cast_8116_wire_constant;
    -- flow-through select operator MUX_8127_inst
    IMA105_8128 <= type_cast_8124_wire_constant when (BITSEL_u8_u1_8122_wire(0) /=  '0') else type_cast_8126_wire_constant;
    -- flow-through select operator MUX_8137_inst
    IMA106_8138 <= type_cast_8134_wire_constant when (BITSEL_u8_u1_8132_wire(0) /=  '0') else type_cast_8136_wire_constant;
    -- flow-through select operator MUX_8147_inst
    IMA107_8148 <= type_cast_8144_wire_constant when (BITSEL_u8_u1_8142_wire(0) /=  '0') else type_cast_8146_wire_constant;
    -- flow-through select operator MUX_8157_inst
    IMA108_8158 <= type_cast_8154_wire_constant when (BITSEL_u8_u1_8152_wire(0) /=  '0') else type_cast_8156_wire_constant;
    -- flow-through select operator MUX_8167_inst
    IMA109_8168 <= type_cast_8164_wire_constant when (BITSEL_u8_u1_8162_wire(0) /=  '0') else type_cast_8166_wire_constant;
    -- flow-through select operator MUX_8177_inst
    IMA110_8178 <= type_cast_8174_wire_constant when (BITSEL_u8_u1_8172_wire(0) /=  '0') else type_cast_8176_wire_constant;
    -- flow-through select operator MUX_8187_inst
    IMA111_8188 <= type_cast_8184_wire_constant when (BITSEL_u8_u1_8182_wire(0) /=  '0') else type_cast_8186_wire_constant;
    -- flow-through select operator MUX_8197_inst
    IMA112_8198 <= type_cast_8194_wire_constant when (BITSEL_u8_u1_8192_wire(0) /=  '0') else type_cast_8196_wire_constant;
    -- flow-through select operator MUX_8207_inst
    IMA113_8208 <= type_cast_8204_wire_constant when (BITSEL_u8_u1_8202_wire(0) /=  '0') else type_cast_8206_wire_constant;
    -- flow-through select operator MUX_8217_inst
    IMA114_8218 <= type_cast_8214_wire_constant when (BITSEL_u8_u1_8212_wire(0) /=  '0') else type_cast_8216_wire_constant;
    -- flow-through select operator MUX_8227_inst
    IMA115_8228 <= type_cast_8224_wire_constant when (BITSEL_u8_u1_8222_wire(0) /=  '0') else type_cast_8226_wire_constant;
    -- flow-through select operator MUX_8237_inst
    IMA116_8238 <= type_cast_8234_wire_constant when (BITSEL_u8_u1_8232_wire(0) /=  '0') else type_cast_8236_wire_constant;
    -- flow-through select operator MUX_8247_inst
    IMA117_8248 <= type_cast_8244_wire_constant when (BITSEL_u8_u1_8242_wire(0) /=  '0') else type_cast_8246_wire_constant;
    -- flow-through select operator MUX_8257_inst
    IMA118_8258 <= type_cast_8254_wire_constant when (BITSEL_u8_u1_8252_wire(0) /=  '0') else type_cast_8256_wire_constant;
    -- flow-through select operator MUX_8267_inst
    IMA119_8268 <= type_cast_8264_wire_constant when (BITSEL_u8_u1_8262_wire(0) /=  '0') else type_cast_8266_wire_constant;
    -- flow-through select operator MUX_8277_inst
    IMA120_8278 <= type_cast_8274_wire_constant when (BITSEL_u8_u1_8272_wire(0) /=  '0') else type_cast_8276_wire_constant;
    -- flow-through select operator MUX_8287_inst
    IMA121_8288 <= type_cast_8284_wire_constant when (BITSEL_u8_u1_8282_wire(0) /=  '0') else type_cast_8286_wire_constant;
    -- flow-through select operator MUX_8297_inst
    IMA122_8298 <= type_cast_8294_wire_constant when (BITSEL_u8_u1_8292_wire(0) /=  '0') else type_cast_8296_wire_constant;
    -- flow-through select operator MUX_8307_inst
    IMA123_8308 <= type_cast_8304_wire_constant when (BITSEL_u8_u1_8302_wire(0) /=  '0') else type_cast_8306_wire_constant;
    -- flow-through select operator MUX_8317_inst
    IMA124_8318 <= type_cast_8314_wire_constant when (BITSEL_u8_u1_8312_wire(0) /=  '0') else type_cast_8316_wire_constant;
    -- flow-through select operator MUX_8327_inst
    IMA125_8328 <= type_cast_8324_wire_constant when (BITSEL_u8_u1_8322_wire(0) /=  '0') else type_cast_8326_wire_constant;
    -- flow-through select operator MUX_8337_inst
    IMA126_8338 <= type_cast_8334_wire_constant when (BITSEL_u8_u1_8332_wire(0) /=  '0') else type_cast_8336_wire_constant;
    -- flow-through select operator MUX_8347_inst
    IMA127_8348 <= type_cast_8344_wire_constant when (BITSEL_u8_u1_8342_wire(0) /=  '0') else type_cast_8346_wire_constant;
    -- flow-through select operator MUX_8355_inst
    IMB0_8356 <= IMA1_7088 when (BITSEL_u8_u1_8352_wire(0) /=  '0') else IMA0_7078;
    -- flow-through select operator MUX_8363_inst
    IMB1_8364 <= IMA3_7108 when (BITSEL_u8_u1_8360_wire(0) /=  '0') else IMA2_7098;
    -- flow-through select operator MUX_8371_inst
    IMB2_8372 <= IMA5_7128 when (BITSEL_u8_u1_8368_wire(0) /=  '0') else IMA4_7118;
    -- flow-through select operator MUX_8379_inst
    IMB3_8380 <= IMA7_7148 when (BITSEL_u8_u1_8376_wire(0) /=  '0') else IMA6_7138;
    -- flow-through select operator MUX_8387_inst
    IMB4_8388 <= IMA9_7168 when (BITSEL_u8_u1_8384_wire(0) /=  '0') else IMA8_7158;
    -- flow-through select operator MUX_8395_inst
    IMB5_8396 <= IMA11_7188 when (BITSEL_u8_u1_8392_wire(0) /=  '0') else IMA10_7178;
    -- flow-through select operator MUX_8403_inst
    IMB6_8404 <= IMA13_7208 when (BITSEL_u8_u1_8400_wire(0) /=  '0') else IMA12_7198;
    -- flow-through select operator MUX_8411_inst
    IMB7_8412 <= IMA15_7228 when (BITSEL_u8_u1_8408_wire(0) /=  '0') else IMA14_7218;
    -- flow-through select operator MUX_8419_inst
    IMB8_8420 <= IMA17_7248 when (BITSEL_u8_u1_8416_wire(0) /=  '0') else IMA16_7238;
    -- flow-through select operator MUX_8427_inst
    IMB9_8428 <= IMA19_7268 when (BITSEL_u8_u1_8424_wire(0) /=  '0') else IMA18_7258;
    -- flow-through select operator MUX_8435_inst
    IMB10_8436 <= IMA21_7288 when (BITSEL_u8_u1_8432_wire(0) /=  '0') else IMA20_7278;
    -- flow-through select operator MUX_8443_inst
    IMB11_8444 <= IMA23_7308 when (BITSEL_u8_u1_8440_wire(0) /=  '0') else IMA22_7298;
    -- flow-through select operator MUX_8451_inst
    IMB12_8452 <= IMA25_7328 when (BITSEL_u8_u1_8448_wire(0) /=  '0') else IMA24_7318;
    -- flow-through select operator MUX_8459_inst
    IMB13_8460 <= IMA27_7348 when (BITSEL_u8_u1_8456_wire(0) /=  '0') else IMA26_7338;
    -- flow-through select operator MUX_8467_inst
    IMB14_8468 <= IMA29_7368 when (BITSEL_u8_u1_8464_wire(0) /=  '0') else IMA28_7358;
    -- flow-through select operator MUX_8475_inst
    IMB15_8476 <= IMA31_7388 when (BITSEL_u8_u1_8472_wire(0) /=  '0') else IMA30_7378;
    -- flow-through select operator MUX_8483_inst
    IMB16_8484 <= IMA33_7408 when (BITSEL_u8_u1_8480_wire(0) /=  '0') else IMA32_7398;
    -- flow-through select operator MUX_8491_inst
    IMB17_8492 <= IMA35_7428 when (BITSEL_u8_u1_8488_wire(0) /=  '0') else IMA34_7418;
    -- flow-through select operator MUX_8499_inst
    IMB18_8500 <= IMA37_7448 when (BITSEL_u8_u1_8496_wire(0) /=  '0') else IMA36_7438;
    -- flow-through select operator MUX_8507_inst
    IMB19_8508 <= IMA39_7468 when (BITSEL_u8_u1_8504_wire(0) /=  '0') else IMA38_7458;
    -- flow-through select operator MUX_8515_inst
    IMB20_8516 <= IMA41_7488 when (BITSEL_u8_u1_8512_wire(0) /=  '0') else IMA40_7478;
    -- flow-through select operator MUX_8523_inst
    IMB21_8524 <= IMA43_7508 when (BITSEL_u8_u1_8520_wire(0) /=  '0') else IMA42_7498;
    -- flow-through select operator MUX_8531_inst
    IMB22_8532 <= IMA45_7528 when (BITSEL_u8_u1_8528_wire(0) /=  '0') else IMA44_7518;
    -- flow-through select operator MUX_8539_inst
    IMB23_8540 <= IMA47_7548 when (BITSEL_u8_u1_8536_wire(0) /=  '0') else IMA46_7538;
    -- flow-through select operator MUX_8547_inst
    IMB24_8548 <= IMA49_7568 when (BITSEL_u8_u1_8544_wire(0) /=  '0') else IMA48_7558;
    -- flow-through select operator MUX_8555_inst
    IMB25_8556 <= IMA51_7588 when (BITSEL_u8_u1_8552_wire(0) /=  '0') else IMA50_7578;
    -- flow-through select operator MUX_8563_inst
    IMB26_8564 <= IMA53_7608 when (BITSEL_u8_u1_8560_wire(0) /=  '0') else IMA52_7598;
    -- flow-through select operator MUX_8571_inst
    IMB27_8572 <= IMA55_7628 when (BITSEL_u8_u1_8568_wire(0) /=  '0') else IMA54_7618;
    -- flow-through select operator MUX_8579_inst
    IMB28_8580 <= IMA57_7648 when (BITSEL_u8_u1_8576_wire(0) /=  '0') else IMA56_7638;
    -- flow-through select operator MUX_8587_inst
    IMB29_8588 <= IMA59_7668 when (BITSEL_u8_u1_8584_wire(0) /=  '0') else IMA58_7658;
    -- flow-through select operator MUX_8595_inst
    IMB30_8596 <= IMA61_7688 when (BITSEL_u8_u1_8592_wire(0) /=  '0') else IMA60_7678;
    -- flow-through select operator MUX_8603_inst
    IMB31_8604 <= IMA63_7708 when (BITSEL_u8_u1_8600_wire(0) /=  '0') else IMA62_7698;
    -- flow-through select operator MUX_8611_inst
    IMB32_8612 <= IMA65_7728 when (BITSEL_u8_u1_8608_wire(0) /=  '0') else IMA64_7718;
    -- flow-through select operator MUX_8619_inst
    IMB33_8620 <= IMA67_7748 when (BITSEL_u8_u1_8616_wire(0) /=  '0') else IMA66_7738;
    -- flow-through select operator MUX_8627_inst
    IMB34_8628 <= IMA69_7768 when (BITSEL_u8_u1_8624_wire(0) /=  '0') else IMA68_7758;
    -- flow-through select operator MUX_8635_inst
    IMB35_8636 <= IMA71_7788 when (BITSEL_u8_u1_8632_wire(0) /=  '0') else IMA70_7778;
    -- flow-through select operator MUX_8643_inst
    IMB36_8644 <= IMA73_7808 when (BITSEL_u8_u1_8640_wire(0) /=  '0') else IMA72_7798;
    -- flow-through select operator MUX_8651_inst
    IMB37_8652 <= IMA75_7828 when (BITSEL_u8_u1_8648_wire(0) /=  '0') else IMA74_7818;
    -- flow-through select operator MUX_8659_inst
    IMB38_8660 <= IMA77_7848 when (BITSEL_u8_u1_8656_wire(0) /=  '0') else IMA76_7838;
    -- flow-through select operator MUX_8667_inst
    IMB39_8668 <= IMA79_7868 when (BITSEL_u8_u1_8664_wire(0) /=  '0') else IMA78_7858;
    -- flow-through select operator MUX_8675_inst
    IMB40_8676 <= IMA81_7888 when (BITSEL_u8_u1_8672_wire(0) /=  '0') else IMA80_7878;
    -- flow-through select operator MUX_8683_inst
    IMB41_8684 <= IMA83_7908 when (BITSEL_u8_u1_8680_wire(0) /=  '0') else IMA82_7898;
    -- flow-through select operator MUX_8691_inst
    IMB42_8692 <= IMA85_7928 when (BITSEL_u8_u1_8688_wire(0) /=  '0') else IMA84_7918;
    -- flow-through select operator MUX_8699_inst
    IMB43_8700 <= IMA87_7948 when (BITSEL_u8_u1_8696_wire(0) /=  '0') else IMA86_7938;
    -- flow-through select operator MUX_8707_inst
    IMB44_8708 <= IMA89_7968 when (BITSEL_u8_u1_8704_wire(0) /=  '0') else IMA88_7958;
    -- flow-through select operator MUX_8715_inst
    IMB45_8716 <= IMA91_7988 when (BITSEL_u8_u1_8712_wire(0) /=  '0') else IMA90_7978;
    -- flow-through select operator MUX_8723_inst
    IMB46_8724 <= IMA93_8008 when (BITSEL_u8_u1_8720_wire(0) /=  '0') else IMA92_7998;
    -- flow-through select operator MUX_8731_inst
    IMB47_8732 <= IMA95_8028 when (BITSEL_u8_u1_8728_wire(0) /=  '0') else IMA94_8018;
    -- flow-through select operator MUX_8739_inst
    IMB48_8740 <= IMA97_8048 when (BITSEL_u8_u1_8736_wire(0) /=  '0') else IMA96_8038;
    -- flow-through select operator MUX_8747_inst
    IMB49_8748 <= IMA99_8068 when (BITSEL_u8_u1_8744_wire(0) /=  '0') else IMA98_8058;
    -- flow-through select operator MUX_8755_inst
    IMB50_8756 <= IMA101_8088 when (BITSEL_u8_u1_8752_wire(0) /=  '0') else IMA100_8078;
    -- flow-through select operator MUX_8763_inst
    IMB51_8764 <= IMA103_8108 when (BITSEL_u8_u1_8760_wire(0) /=  '0') else IMA102_8098;
    -- flow-through select operator MUX_8771_inst
    IMB52_8772 <= IMA105_8128 when (BITSEL_u8_u1_8768_wire(0) /=  '0') else IMA104_8118;
    -- flow-through select operator MUX_8779_inst
    IMB53_8780 <= IMA107_8148 when (BITSEL_u8_u1_8776_wire(0) /=  '0') else IMA106_8138;
    -- flow-through select operator MUX_8787_inst
    IMB54_8788 <= IMA109_8168 when (BITSEL_u8_u1_8784_wire(0) /=  '0') else IMA108_8158;
    -- flow-through select operator MUX_8795_inst
    IMB55_8796 <= IMA111_8188 when (BITSEL_u8_u1_8792_wire(0) /=  '0') else IMA110_8178;
    -- flow-through select operator MUX_8803_inst
    IMB56_8804 <= IMA113_8208 when (BITSEL_u8_u1_8800_wire(0) /=  '0') else IMA112_8198;
    -- flow-through select operator MUX_8811_inst
    IMB57_8812 <= IMA115_8228 when (BITSEL_u8_u1_8808_wire(0) /=  '0') else IMA114_8218;
    -- flow-through select operator MUX_8819_inst
    IMB58_8820 <= IMA117_8248 when (BITSEL_u8_u1_8816_wire(0) /=  '0') else IMA116_8238;
    -- flow-through select operator MUX_8827_inst
    IMB59_8828 <= IMA119_8268 when (BITSEL_u8_u1_8824_wire(0) /=  '0') else IMA118_8258;
    -- flow-through select operator MUX_8835_inst
    IMB60_8836 <= IMA121_8288 when (BITSEL_u8_u1_8832_wire(0) /=  '0') else IMA120_8278;
    -- flow-through select operator MUX_8843_inst
    IMB61_8844 <= IMA123_8308 when (BITSEL_u8_u1_8840_wire(0) /=  '0') else IMA122_8298;
    -- flow-through select operator MUX_8851_inst
    IMB62_8852 <= IMA125_8328 when (BITSEL_u8_u1_8848_wire(0) /=  '0') else IMA124_8318;
    -- flow-through select operator MUX_8859_inst
    IMB63_8860 <= IMA127_8348 when (BITSEL_u8_u1_8856_wire(0) /=  '0') else IMA126_8338;
    -- flow-through select operator MUX_8867_inst
    IMC0_8868 <= IMB1_8364 when (BITSEL_u8_u1_8864_wire(0) /=  '0') else IMB0_8356;
    -- flow-through select operator MUX_8875_inst
    IMC1_8876 <= IMB3_8380 when (BITSEL_u8_u1_8872_wire(0) /=  '0') else IMB2_8372;
    -- flow-through select operator MUX_8883_inst
    IMC2_8884 <= IMB5_8396 when (BITSEL_u8_u1_8880_wire(0) /=  '0') else IMB4_8388;
    -- flow-through select operator MUX_8891_inst
    IMC3_8892 <= IMB7_8412 when (BITSEL_u8_u1_8888_wire(0) /=  '0') else IMB6_8404;
    -- flow-through select operator MUX_8899_inst
    IMC4_8900 <= IMB9_8428 when (BITSEL_u8_u1_8896_wire(0) /=  '0') else IMB8_8420;
    -- flow-through select operator MUX_8907_inst
    IMC5_8908 <= IMB11_8444 when (BITSEL_u8_u1_8904_wire(0) /=  '0') else IMB10_8436;
    -- flow-through select operator MUX_8915_inst
    IMC6_8916 <= IMB13_8460 when (BITSEL_u8_u1_8912_wire(0) /=  '0') else IMB12_8452;
    -- flow-through select operator MUX_8923_inst
    IMC7_8924 <= IMB15_8476 when (BITSEL_u8_u1_8920_wire(0) /=  '0') else IMB14_8468;
    -- flow-through select operator MUX_8931_inst
    IMC8_8932 <= IMB17_8492 when (BITSEL_u8_u1_8928_wire(0) /=  '0') else IMB16_8484;
    -- flow-through select operator MUX_8939_inst
    IMC9_8940 <= IMB19_8508 when (BITSEL_u8_u1_8936_wire(0) /=  '0') else IMB18_8500;
    -- flow-through select operator MUX_8947_inst
    IMC10_8948 <= IMB21_8524 when (BITSEL_u8_u1_8944_wire(0) /=  '0') else IMB20_8516;
    -- flow-through select operator MUX_8955_inst
    IMC11_8956 <= IMB23_8540 when (BITSEL_u8_u1_8952_wire(0) /=  '0') else IMB22_8532;
    -- flow-through select operator MUX_8963_inst
    IMC12_8964 <= IMB25_8556 when (BITSEL_u8_u1_8960_wire(0) /=  '0') else IMB24_8548;
    -- flow-through select operator MUX_8971_inst
    IMC13_8972 <= IMB27_8572 when (BITSEL_u8_u1_8968_wire(0) /=  '0') else IMB26_8564;
    -- flow-through select operator MUX_8979_inst
    IMC14_8980 <= IMB29_8588 when (BITSEL_u8_u1_8976_wire(0) /=  '0') else IMB28_8580;
    -- flow-through select operator MUX_8987_inst
    IMC15_8988 <= IMB31_8604 when (BITSEL_u8_u1_8984_wire(0) /=  '0') else IMB30_8596;
    -- flow-through select operator MUX_8995_inst
    IMC16_8996 <= IMB33_8620 when (BITSEL_u8_u1_8992_wire(0) /=  '0') else IMB32_8612;
    -- flow-through select operator MUX_9003_inst
    IMC17_9004 <= IMB35_8636 when (BITSEL_u8_u1_9000_wire(0) /=  '0') else IMB34_8628;
    -- flow-through select operator MUX_9011_inst
    IMC18_9012 <= IMB37_8652 when (BITSEL_u8_u1_9008_wire(0) /=  '0') else IMB36_8644;
    -- flow-through select operator MUX_9019_inst
    IMC19_9020 <= IMB39_8668 when (BITSEL_u8_u1_9016_wire(0) /=  '0') else IMB38_8660;
    -- flow-through select operator MUX_9027_inst
    IMC20_9028 <= IMB41_8684 when (BITSEL_u8_u1_9024_wire(0) /=  '0') else IMB40_8676;
    -- flow-through select operator MUX_9035_inst
    IMC21_9036 <= IMB43_8700 when (BITSEL_u8_u1_9032_wire(0) /=  '0') else IMB42_8692;
    -- flow-through select operator MUX_9043_inst
    IMC22_9044 <= IMB45_8716 when (BITSEL_u8_u1_9040_wire(0) /=  '0') else IMB44_8708;
    -- flow-through select operator MUX_9051_inst
    IMC23_9052 <= IMB47_8732 when (BITSEL_u8_u1_9048_wire(0) /=  '0') else IMB46_8724;
    -- flow-through select operator MUX_9059_inst
    IMC24_9060 <= IMB49_8748 when (BITSEL_u8_u1_9056_wire(0) /=  '0') else IMB48_8740;
    -- flow-through select operator MUX_9067_inst
    IMC25_9068 <= IMB51_8764 when (BITSEL_u8_u1_9064_wire(0) /=  '0') else IMB50_8756;
    -- flow-through select operator MUX_9075_inst
    IMC26_9076 <= IMB53_8780 when (BITSEL_u8_u1_9072_wire(0) /=  '0') else IMB52_8772;
    -- flow-through select operator MUX_9083_inst
    IMC27_9084 <= IMB55_8796 when (BITSEL_u8_u1_9080_wire(0) /=  '0') else IMB54_8788;
    -- flow-through select operator MUX_9091_inst
    IMC28_9092 <= IMB57_8812 when (BITSEL_u8_u1_9088_wire(0) /=  '0') else IMB56_8804;
    -- flow-through select operator MUX_9099_inst
    IMC29_9100 <= IMB59_8828 when (BITSEL_u8_u1_9096_wire(0) /=  '0') else IMB58_8820;
    -- flow-through select operator MUX_9107_inst
    IMC30_9108 <= IMB61_8844 when (BITSEL_u8_u1_9104_wire(0) /=  '0') else IMB60_8836;
    -- flow-through select operator MUX_9115_inst
    IMC31_9116 <= IMB63_8860 when (BITSEL_u8_u1_9112_wire(0) /=  '0') else IMB62_8852;
    -- flow-through select operator MUX_9123_inst
    IMD0_9124 <= IMC1_8876 when (BITSEL_u8_u1_9120_wire(0) /=  '0') else IMC0_8868;
    -- flow-through select operator MUX_9131_inst
    IMD1_9132 <= IMC3_8892 when (BITSEL_u8_u1_9128_wire(0) /=  '0') else IMC2_8884;
    -- flow-through select operator MUX_9139_inst
    IMD2_9140 <= IMC5_8908 when (BITSEL_u8_u1_9136_wire(0) /=  '0') else IMC4_8900;
    -- flow-through select operator MUX_9147_inst
    IMD3_9148 <= IMC7_8924 when (BITSEL_u8_u1_9144_wire(0) /=  '0') else IMC6_8916;
    -- flow-through select operator MUX_9155_inst
    IMD4_9156 <= IMC9_8940 when (BITSEL_u8_u1_9152_wire(0) /=  '0') else IMC8_8932;
    -- flow-through select operator MUX_9163_inst
    IMD5_9164 <= IMC11_8956 when (BITSEL_u8_u1_9160_wire(0) /=  '0') else IMC10_8948;
    -- flow-through select operator MUX_9171_inst
    IMD6_9172 <= IMC13_8972 when (BITSEL_u8_u1_9168_wire(0) /=  '0') else IMC12_8964;
    -- flow-through select operator MUX_9179_inst
    IMD7_9180 <= IMC15_8988 when (BITSEL_u8_u1_9176_wire(0) /=  '0') else IMC14_8980;
    -- flow-through select operator MUX_9187_inst
    IMD8_9188 <= IMC17_9004 when (BITSEL_u8_u1_9184_wire(0) /=  '0') else IMC16_8996;
    -- flow-through select operator MUX_9195_inst
    IMD9_9196 <= IMC19_9020 when (BITSEL_u8_u1_9192_wire(0) /=  '0') else IMC18_9012;
    -- flow-through select operator MUX_9203_inst
    IMD10_9204 <= IMC21_9036 when (BITSEL_u8_u1_9200_wire(0) /=  '0') else IMC20_9028;
    -- flow-through select operator MUX_9211_inst
    IMD11_9212 <= IMC23_9052 when (BITSEL_u8_u1_9208_wire(0) /=  '0') else IMC22_9044;
    -- flow-through select operator MUX_9219_inst
    IMD12_9220 <= IMC25_9068 when (BITSEL_u8_u1_9216_wire(0) /=  '0') else IMC24_9060;
    -- flow-through select operator MUX_9227_inst
    IMD13_9228 <= IMC27_9084 when (BITSEL_u8_u1_9224_wire(0) /=  '0') else IMC26_9076;
    -- flow-through select operator MUX_9235_inst
    IMD14_9236 <= IMC29_9100 when (BITSEL_u8_u1_9232_wire(0) /=  '0') else IMC28_9092;
    -- flow-through select operator MUX_9243_inst
    IMD15_9244 <= IMC31_9116 when (BITSEL_u8_u1_9240_wire(0) /=  '0') else IMC30_9108;
    -- flow-through select operator MUX_9251_inst
    IME0_9252 <= IMD1_9132 when (BITSEL_u8_u1_9248_wire(0) /=  '0') else IMD0_9124;
    -- flow-through select operator MUX_9259_inst
    IME1_9260 <= IMD3_9148 when (BITSEL_u8_u1_9256_wire(0) /=  '0') else IMD2_9140;
    -- flow-through select operator MUX_9267_inst
    IME2_9268 <= IMD5_9164 when (BITSEL_u8_u1_9264_wire(0) /=  '0') else IMD4_9156;
    -- flow-through select operator MUX_9275_inst
    IME3_9276 <= IMD7_9180 when (BITSEL_u8_u1_9272_wire(0) /=  '0') else IMD6_9172;
    -- flow-through select operator MUX_9283_inst
    IME4_9284 <= IMD9_9196 when (BITSEL_u8_u1_9280_wire(0) /=  '0') else IMD8_9188;
    -- flow-through select operator MUX_9291_inst
    IME5_9292 <= IMD11_9212 when (BITSEL_u8_u1_9288_wire(0) /=  '0') else IMD10_9204;
    -- flow-through select operator MUX_9299_inst
    IME6_9300 <= IMD13_9228 when (BITSEL_u8_u1_9296_wire(0) /=  '0') else IMD12_9220;
    -- flow-through select operator MUX_9307_inst
    IME7_9308 <= IMD15_9244 when (BITSEL_u8_u1_9304_wire(0) /=  '0') else IMD14_9236;
    -- flow-through select operator MUX_9315_inst
    IMF0_9316 <= IME1_9260 when (BITSEL_u8_u1_9312_wire(0) /=  '0') else IME0_9252;
    -- flow-through select operator MUX_9323_inst
    IMF1_9324 <= IME3_9276 when (BITSEL_u8_u1_9320_wire(0) /=  '0') else IME2_9268;
    -- flow-through select operator MUX_9331_inst
    IMF2_9332 <= IME5_9292 when (BITSEL_u8_u1_9328_wire(0) /=  '0') else IME4_9284;
    -- flow-through select operator MUX_9339_inst
    IMF3_9340 <= IME7_9308 when (BITSEL_u8_u1_9336_wire(0) /=  '0') else IME6_9300;
    -- flow-through select operator MUX_9347_inst
    IMG0_9348 <= IMF1_9324 when (BITSEL_u8_u1_9344_wire(0) /=  '0') else IMF0_9316;
    -- flow-through select operator MUX_9355_inst
    IMG1_9356 <= IMF3_9340 when (BITSEL_u8_u1_9352_wire(0) /=  '0') else IMF2_9332;
    -- flow-through select operator MUX_9363_inst
    s_out_buffer <= IMG1_9356 when (BITSEL_u8_u1_9360_wire(0) /=  '0') else IMG0_9348;
    -- binary operator BITSEL_u8_u1_7072_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7071_wire_constant, tmp_var);
      BITSEL_u8_u1_7072_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_7082_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7081_wire_constant, tmp_var);
      BITSEL_u8_u1_7082_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_7092_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7091_wire_constant, tmp_var);
      BITSEL_u8_u1_7092_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_7102_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7101_wire_constant, tmp_var);
      BITSEL_u8_u1_7102_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_7112_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7111_wire_constant, tmp_var);
      BITSEL_u8_u1_7112_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_7122_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7121_wire_constant, tmp_var);
      BITSEL_u8_u1_7122_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_7132_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7131_wire_constant, tmp_var);
      BITSEL_u8_u1_7132_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_7142_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7141_wire_constant, tmp_var);
      BITSEL_u8_u1_7142_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_7152_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7151_wire_constant, tmp_var);
      BITSEL_u8_u1_7152_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_7162_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7161_wire_constant, tmp_var);
      BITSEL_u8_u1_7162_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_7172_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7171_wire_constant, tmp_var);
      BITSEL_u8_u1_7172_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_7182_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7181_wire_constant, tmp_var);
      BITSEL_u8_u1_7182_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_7192_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7191_wire_constant, tmp_var);
      BITSEL_u8_u1_7192_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_7202_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7201_wire_constant, tmp_var);
      BITSEL_u8_u1_7202_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_7212_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7211_wire_constant, tmp_var);
      BITSEL_u8_u1_7212_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_7222_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7221_wire_constant, tmp_var);
      BITSEL_u8_u1_7222_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_7232_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7231_wire_constant, tmp_var);
      BITSEL_u8_u1_7232_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_7242_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7241_wire_constant, tmp_var);
      BITSEL_u8_u1_7242_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_7252_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7251_wire_constant, tmp_var);
      BITSEL_u8_u1_7252_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_7262_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7261_wire_constant, tmp_var);
      BITSEL_u8_u1_7262_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_7272_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7271_wire_constant, tmp_var);
      BITSEL_u8_u1_7272_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_7282_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7281_wire_constant, tmp_var);
      BITSEL_u8_u1_7282_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_7292_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7291_wire_constant, tmp_var);
      BITSEL_u8_u1_7292_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_7302_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7301_wire_constant, tmp_var);
      BITSEL_u8_u1_7302_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_7312_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7311_wire_constant, tmp_var);
      BITSEL_u8_u1_7312_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_7322_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7321_wire_constant, tmp_var);
      BITSEL_u8_u1_7322_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_7332_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7331_wire_constant, tmp_var);
      BITSEL_u8_u1_7332_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_7342_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7341_wire_constant, tmp_var);
      BITSEL_u8_u1_7342_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_7352_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7351_wire_constant, tmp_var);
      BITSEL_u8_u1_7352_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_7362_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7361_wire_constant, tmp_var);
      BITSEL_u8_u1_7362_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_7372_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7371_wire_constant, tmp_var);
      BITSEL_u8_u1_7372_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_7382_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7381_wire_constant, tmp_var);
      BITSEL_u8_u1_7382_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_7392_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7391_wire_constant, tmp_var);
      BITSEL_u8_u1_7392_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_7402_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7401_wire_constant, tmp_var);
      BITSEL_u8_u1_7402_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_7412_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7411_wire_constant, tmp_var);
      BITSEL_u8_u1_7412_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_7422_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7421_wire_constant, tmp_var);
      BITSEL_u8_u1_7422_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_7432_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7431_wire_constant, tmp_var);
      BITSEL_u8_u1_7432_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_7442_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7441_wire_constant, tmp_var);
      BITSEL_u8_u1_7442_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_7452_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7451_wire_constant, tmp_var);
      BITSEL_u8_u1_7452_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_7462_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7461_wire_constant, tmp_var);
      BITSEL_u8_u1_7462_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_7472_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7471_wire_constant, tmp_var);
      BITSEL_u8_u1_7472_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_7482_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7481_wire_constant, tmp_var);
      BITSEL_u8_u1_7482_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_7492_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7491_wire_constant, tmp_var);
      BITSEL_u8_u1_7492_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_7502_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7501_wire_constant, tmp_var);
      BITSEL_u8_u1_7502_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_7512_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7511_wire_constant, tmp_var);
      BITSEL_u8_u1_7512_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_7522_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7521_wire_constant, tmp_var);
      BITSEL_u8_u1_7522_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_7532_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7531_wire_constant, tmp_var);
      BITSEL_u8_u1_7532_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_7542_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7541_wire_constant, tmp_var);
      BITSEL_u8_u1_7542_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_7552_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7551_wire_constant, tmp_var);
      BITSEL_u8_u1_7552_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_7562_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7561_wire_constant, tmp_var);
      BITSEL_u8_u1_7562_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_7572_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7571_wire_constant, tmp_var);
      BITSEL_u8_u1_7572_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_7582_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7581_wire_constant, tmp_var);
      BITSEL_u8_u1_7582_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_7592_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7591_wire_constant, tmp_var);
      BITSEL_u8_u1_7592_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_7602_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7601_wire_constant, tmp_var);
      BITSEL_u8_u1_7602_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_7612_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7611_wire_constant, tmp_var);
      BITSEL_u8_u1_7612_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_7622_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7621_wire_constant, tmp_var);
      BITSEL_u8_u1_7622_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_7632_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7631_wire_constant, tmp_var);
      BITSEL_u8_u1_7632_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_7642_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7641_wire_constant, tmp_var);
      BITSEL_u8_u1_7642_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_7652_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7651_wire_constant, tmp_var);
      BITSEL_u8_u1_7652_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_7662_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7661_wire_constant, tmp_var);
      BITSEL_u8_u1_7662_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_7672_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7671_wire_constant, tmp_var);
      BITSEL_u8_u1_7672_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_7682_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7681_wire_constant, tmp_var);
      BITSEL_u8_u1_7682_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_7692_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7691_wire_constant, tmp_var);
      BITSEL_u8_u1_7692_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_7702_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7701_wire_constant, tmp_var);
      BITSEL_u8_u1_7702_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_7712_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7711_wire_constant, tmp_var);
      BITSEL_u8_u1_7712_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_7722_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7721_wire_constant, tmp_var);
      BITSEL_u8_u1_7722_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_7732_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7731_wire_constant, tmp_var);
      BITSEL_u8_u1_7732_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_7742_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7741_wire_constant, tmp_var);
      BITSEL_u8_u1_7742_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_7752_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7751_wire_constant, tmp_var);
      BITSEL_u8_u1_7752_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_7762_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7761_wire_constant, tmp_var);
      BITSEL_u8_u1_7762_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_7772_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7771_wire_constant, tmp_var);
      BITSEL_u8_u1_7772_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_7782_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7781_wire_constant, tmp_var);
      BITSEL_u8_u1_7782_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_7792_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7791_wire_constant, tmp_var);
      BITSEL_u8_u1_7792_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_7802_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7801_wire_constant, tmp_var);
      BITSEL_u8_u1_7802_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_7812_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7811_wire_constant, tmp_var);
      BITSEL_u8_u1_7812_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_7822_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7821_wire_constant, tmp_var);
      BITSEL_u8_u1_7822_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_7832_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7831_wire_constant, tmp_var);
      BITSEL_u8_u1_7832_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_7842_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7841_wire_constant, tmp_var);
      BITSEL_u8_u1_7842_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_7852_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7851_wire_constant, tmp_var);
      BITSEL_u8_u1_7852_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_7862_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7861_wire_constant, tmp_var);
      BITSEL_u8_u1_7862_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_7872_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7871_wire_constant, tmp_var);
      BITSEL_u8_u1_7872_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_7882_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7881_wire_constant, tmp_var);
      BITSEL_u8_u1_7882_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_7892_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7891_wire_constant, tmp_var);
      BITSEL_u8_u1_7892_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_7902_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7901_wire_constant, tmp_var);
      BITSEL_u8_u1_7902_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_7912_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7911_wire_constant, tmp_var);
      BITSEL_u8_u1_7912_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_7922_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7921_wire_constant, tmp_var);
      BITSEL_u8_u1_7922_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_7932_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7931_wire_constant, tmp_var);
      BITSEL_u8_u1_7932_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_7942_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7941_wire_constant, tmp_var);
      BITSEL_u8_u1_7942_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_7952_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7951_wire_constant, tmp_var);
      BITSEL_u8_u1_7952_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_7962_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7961_wire_constant, tmp_var);
      BITSEL_u8_u1_7962_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_7972_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7971_wire_constant, tmp_var);
      BITSEL_u8_u1_7972_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_7982_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7981_wire_constant, tmp_var);
      BITSEL_u8_u1_7982_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_7992_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_7991_wire_constant, tmp_var);
      BITSEL_u8_u1_7992_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8002_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8001_wire_constant, tmp_var);
      BITSEL_u8_u1_8002_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8012_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8011_wire_constant, tmp_var);
      BITSEL_u8_u1_8012_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8022_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8021_wire_constant, tmp_var);
      BITSEL_u8_u1_8022_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8032_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8031_wire_constant, tmp_var);
      BITSEL_u8_u1_8032_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8042_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8041_wire_constant, tmp_var);
      BITSEL_u8_u1_8042_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8052_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8051_wire_constant, tmp_var);
      BITSEL_u8_u1_8052_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8062_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8061_wire_constant, tmp_var);
      BITSEL_u8_u1_8062_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8072_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8071_wire_constant, tmp_var);
      BITSEL_u8_u1_8072_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8082_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8081_wire_constant, tmp_var);
      BITSEL_u8_u1_8082_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8092_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8091_wire_constant, tmp_var);
      BITSEL_u8_u1_8092_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8102_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8101_wire_constant, tmp_var);
      BITSEL_u8_u1_8102_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8112_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8111_wire_constant, tmp_var);
      BITSEL_u8_u1_8112_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8122_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8121_wire_constant, tmp_var);
      BITSEL_u8_u1_8122_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8132_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8131_wire_constant, tmp_var);
      BITSEL_u8_u1_8132_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8142_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8141_wire_constant, tmp_var);
      BITSEL_u8_u1_8142_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8152_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8151_wire_constant, tmp_var);
      BITSEL_u8_u1_8152_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8162_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8161_wire_constant, tmp_var);
      BITSEL_u8_u1_8162_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8172_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8171_wire_constant, tmp_var);
      BITSEL_u8_u1_8172_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8182_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8181_wire_constant, tmp_var);
      BITSEL_u8_u1_8182_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8192_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8191_wire_constant, tmp_var);
      BITSEL_u8_u1_8192_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8202_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8201_wire_constant, tmp_var);
      BITSEL_u8_u1_8202_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8212_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8211_wire_constant, tmp_var);
      BITSEL_u8_u1_8212_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8222_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8221_wire_constant, tmp_var);
      BITSEL_u8_u1_8222_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8232_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8231_wire_constant, tmp_var);
      BITSEL_u8_u1_8232_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8242_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8241_wire_constant, tmp_var);
      BITSEL_u8_u1_8242_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8252_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8251_wire_constant, tmp_var);
      BITSEL_u8_u1_8252_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8262_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8261_wire_constant, tmp_var);
      BITSEL_u8_u1_8262_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8272_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8271_wire_constant, tmp_var);
      BITSEL_u8_u1_8272_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8282_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8281_wire_constant, tmp_var);
      BITSEL_u8_u1_8282_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8292_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8291_wire_constant, tmp_var);
      BITSEL_u8_u1_8292_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8302_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8301_wire_constant, tmp_var);
      BITSEL_u8_u1_8302_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8312_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8311_wire_constant, tmp_var);
      BITSEL_u8_u1_8312_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8322_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8321_wire_constant, tmp_var);
      BITSEL_u8_u1_8322_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8332_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8331_wire_constant, tmp_var);
      BITSEL_u8_u1_8332_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8342_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8341_wire_constant, tmp_var);
      BITSEL_u8_u1_8342_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8352_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8351_wire_constant, tmp_var);
      BITSEL_u8_u1_8352_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8360_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8359_wire_constant, tmp_var);
      BITSEL_u8_u1_8360_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8368_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8367_wire_constant, tmp_var);
      BITSEL_u8_u1_8368_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8376_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8375_wire_constant, tmp_var);
      BITSEL_u8_u1_8376_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8384_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8383_wire_constant, tmp_var);
      BITSEL_u8_u1_8384_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8392_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8391_wire_constant, tmp_var);
      BITSEL_u8_u1_8392_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8400_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8399_wire_constant, tmp_var);
      BITSEL_u8_u1_8400_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8408_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8407_wire_constant, tmp_var);
      BITSEL_u8_u1_8408_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8416_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8415_wire_constant, tmp_var);
      BITSEL_u8_u1_8416_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8424_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8423_wire_constant, tmp_var);
      BITSEL_u8_u1_8424_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8432_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8431_wire_constant, tmp_var);
      BITSEL_u8_u1_8432_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8440_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8439_wire_constant, tmp_var);
      BITSEL_u8_u1_8440_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8448_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8447_wire_constant, tmp_var);
      BITSEL_u8_u1_8448_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8456_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8455_wire_constant, tmp_var);
      BITSEL_u8_u1_8456_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8464_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8463_wire_constant, tmp_var);
      BITSEL_u8_u1_8464_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8472_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8471_wire_constant, tmp_var);
      BITSEL_u8_u1_8472_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8480_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8479_wire_constant, tmp_var);
      BITSEL_u8_u1_8480_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8488_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8487_wire_constant, tmp_var);
      BITSEL_u8_u1_8488_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8496_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8495_wire_constant, tmp_var);
      BITSEL_u8_u1_8496_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8504_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8503_wire_constant, tmp_var);
      BITSEL_u8_u1_8504_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8512_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8511_wire_constant, tmp_var);
      BITSEL_u8_u1_8512_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8520_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8519_wire_constant, tmp_var);
      BITSEL_u8_u1_8520_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8528_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8527_wire_constant, tmp_var);
      BITSEL_u8_u1_8528_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8536_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8535_wire_constant, tmp_var);
      BITSEL_u8_u1_8536_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8544_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8543_wire_constant, tmp_var);
      BITSEL_u8_u1_8544_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8552_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8551_wire_constant, tmp_var);
      BITSEL_u8_u1_8552_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8560_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8559_wire_constant, tmp_var);
      BITSEL_u8_u1_8560_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8568_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8567_wire_constant, tmp_var);
      BITSEL_u8_u1_8568_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8576_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8575_wire_constant, tmp_var);
      BITSEL_u8_u1_8576_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8584_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8583_wire_constant, tmp_var);
      BITSEL_u8_u1_8584_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8592_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8591_wire_constant, tmp_var);
      BITSEL_u8_u1_8592_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8600_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8599_wire_constant, tmp_var);
      BITSEL_u8_u1_8600_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8608_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8607_wire_constant, tmp_var);
      BITSEL_u8_u1_8608_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8616_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8615_wire_constant, tmp_var);
      BITSEL_u8_u1_8616_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8624_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8623_wire_constant, tmp_var);
      BITSEL_u8_u1_8624_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8632_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8631_wire_constant, tmp_var);
      BITSEL_u8_u1_8632_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8640_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8639_wire_constant, tmp_var);
      BITSEL_u8_u1_8640_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8648_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8647_wire_constant, tmp_var);
      BITSEL_u8_u1_8648_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8656_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8655_wire_constant, tmp_var);
      BITSEL_u8_u1_8656_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8664_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8663_wire_constant, tmp_var);
      BITSEL_u8_u1_8664_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8672_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8671_wire_constant, tmp_var);
      BITSEL_u8_u1_8672_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8680_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8679_wire_constant, tmp_var);
      BITSEL_u8_u1_8680_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8688_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8687_wire_constant, tmp_var);
      BITSEL_u8_u1_8688_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8696_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8695_wire_constant, tmp_var);
      BITSEL_u8_u1_8696_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8704_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8703_wire_constant, tmp_var);
      BITSEL_u8_u1_8704_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8712_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8711_wire_constant, tmp_var);
      BITSEL_u8_u1_8712_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8720_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8719_wire_constant, tmp_var);
      BITSEL_u8_u1_8720_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8728_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8727_wire_constant, tmp_var);
      BITSEL_u8_u1_8728_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8736_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8735_wire_constant, tmp_var);
      BITSEL_u8_u1_8736_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8744_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8743_wire_constant, tmp_var);
      BITSEL_u8_u1_8744_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8752_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8751_wire_constant, tmp_var);
      BITSEL_u8_u1_8752_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8760_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8759_wire_constant, tmp_var);
      BITSEL_u8_u1_8760_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8768_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8767_wire_constant, tmp_var);
      BITSEL_u8_u1_8768_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8776_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8775_wire_constant, tmp_var);
      BITSEL_u8_u1_8776_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8784_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8783_wire_constant, tmp_var);
      BITSEL_u8_u1_8784_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8792_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8791_wire_constant, tmp_var);
      BITSEL_u8_u1_8792_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8800_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8799_wire_constant, tmp_var);
      BITSEL_u8_u1_8800_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8808_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8807_wire_constant, tmp_var);
      BITSEL_u8_u1_8808_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8816_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8815_wire_constant, tmp_var);
      BITSEL_u8_u1_8816_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8824_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8823_wire_constant, tmp_var);
      BITSEL_u8_u1_8824_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8832_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8831_wire_constant, tmp_var);
      BITSEL_u8_u1_8832_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8840_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8839_wire_constant, tmp_var);
      BITSEL_u8_u1_8840_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8848_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8847_wire_constant, tmp_var);
      BITSEL_u8_u1_8848_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8856_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8855_wire_constant, tmp_var);
      BITSEL_u8_u1_8856_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8864_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8863_wire_constant, tmp_var);
      BITSEL_u8_u1_8864_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8872_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8871_wire_constant, tmp_var);
      BITSEL_u8_u1_8872_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8880_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8879_wire_constant, tmp_var);
      BITSEL_u8_u1_8880_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8888_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8887_wire_constant, tmp_var);
      BITSEL_u8_u1_8888_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8896_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8895_wire_constant, tmp_var);
      BITSEL_u8_u1_8896_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8904_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8903_wire_constant, tmp_var);
      BITSEL_u8_u1_8904_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8912_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8911_wire_constant, tmp_var);
      BITSEL_u8_u1_8912_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8920_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8919_wire_constant, tmp_var);
      BITSEL_u8_u1_8920_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8928_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8927_wire_constant, tmp_var);
      BITSEL_u8_u1_8928_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8936_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8935_wire_constant, tmp_var);
      BITSEL_u8_u1_8936_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8944_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8943_wire_constant, tmp_var);
      BITSEL_u8_u1_8944_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8952_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8951_wire_constant, tmp_var);
      BITSEL_u8_u1_8952_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8960_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8959_wire_constant, tmp_var);
      BITSEL_u8_u1_8960_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8968_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8967_wire_constant, tmp_var);
      BITSEL_u8_u1_8968_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8976_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8975_wire_constant, tmp_var);
      BITSEL_u8_u1_8976_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8984_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8983_wire_constant, tmp_var);
      BITSEL_u8_u1_8984_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_8992_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8991_wire_constant, tmp_var);
      BITSEL_u8_u1_8992_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_9000_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_8999_wire_constant, tmp_var);
      BITSEL_u8_u1_9000_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_9008_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_9007_wire_constant, tmp_var);
      BITSEL_u8_u1_9008_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_9016_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_9015_wire_constant, tmp_var);
      BITSEL_u8_u1_9016_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_9024_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_9023_wire_constant, tmp_var);
      BITSEL_u8_u1_9024_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_9032_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_9031_wire_constant, tmp_var);
      BITSEL_u8_u1_9032_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_9040_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_9039_wire_constant, tmp_var);
      BITSEL_u8_u1_9040_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_9048_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_9047_wire_constant, tmp_var);
      BITSEL_u8_u1_9048_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_9056_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_9055_wire_constant, tmp_var);
      BITSEL_u8_u1_9056_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_9064_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_9063_wire_constant, tmp_var);
      BITSEL_u8_u1_9064_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_9072_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_9071_wire_constant, tmp_var);
      BITSEL_u8_u1_9072_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_9080_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_9079_wire_constant, tmp_var);
      BITSEL_u8_u1_9080_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_9088_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_9087_wire_constant, tmp_var);
      BITSEL_u8_u1_9088_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_9096_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_9095_wire_constant, tmp_var);
      BITSEL_u8_u1_9096_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_9104_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_9103_wire_constant, tmp_var);
      BITSEL_u8_u1_9104_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_9112_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_9111_wire_constant, tmp_var);
      BITSEL_u8_u1_9112_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_9120_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_9119_wire_constant, tmp_var);
      BITSEL_u8_u1_9120_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_9128_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_9127_wire_constant, tmp_var);
      BITSEL_u8_u1_9128_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_9136_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_9135_wire_constant, tmp_var);
      BITSEL_u8_u1_9136_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_9144_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_9143_wire_constant, tmp_var);
      BITSEL_u8_u1_9144_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_9152_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_9151_wire_constant, tmp_var);
      BITSEL_u8_u1_9152_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_9160_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_9159_wire_constant, tmp_var);
      BITSEL_u8_u1_9160_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_9168_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_9167_wire_constant, tmp_var);
      BITSEL_u8_u1_9168_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_9176_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_9175_wire_constant, tmp_var);
      BITSEL_u8_u1_9176_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_9184_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_9183_wire_constant, tmp_var);
      BITSEL_u8_u1_9184_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_9192_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_9191_wire_constant, tmp_var);
      BITSEL_u8_u1_9192_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_9200_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_9199_wire_constant, tmp_var);
      BITSEL_u8_u1_9200_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_9208_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_9207_wire_constant, tmp_var);
      BITSEL_u8_u1_9208_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_9216_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_9215_wire_constant, tmp_var);
      BITSEL_u8_u1_9216_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_9224_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_9223_wire_constant, tmp_var);
      BITSEL_u8_u1_9224_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_9232_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_9231_wire_constant, tmp_var);
      BITSEL_u8_u1_9232_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_9240_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_9239_wire_constant, tmp_var);
      BITSEL_u8_u1_9240_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_9248_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_9247_wire_constant, tmp_var);
      BITSEL_u8_u1_9248_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_9256_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_9255_wire_constant, tmp_var);
      BITSEL_u8_u1_9256_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_9264_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_9263_wire_constant, tmp_var);
      BITSEL_u8_u1_9264_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_9272_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_9271_wire_constant, tmp_var);
      BITSEL_u8_u1_9272_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_9280_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_9279_wire_constant, tmp_var);
      BITSEL_u8_u1_9280_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_9288_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_9287_wire_constant, tmp_var);
      BITSEL_u8_u1_9288_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_9296_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_9295_wire_constant, tmp_var);
      BITSEL_u8_u1_9296_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_9304_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_9303_wire_constant, tmp_var);
      BITSEL_u8_u1_9304_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_9312_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_9311_wire_constant, tmp_var);
      BITSEL_u8_u1_9312_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_9320_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_9319_wire_constant, tmp_var);
      BITSEL_u8_u1_9320_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_9328_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_9327_wire_constant, tmp_var);
      BITSEL_u8_u1_9328_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_9336_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_9335_wire_constant, tmp_var);
      BITSEL_u8_u1_9336_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_9344_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_9343_wire_constant, tmp_var);
      BITSEL_u8_u1_9344_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_9352_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_9351_wire_constant, tmp_var);
      BITSEL_u8_u1_9352_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_9360_inst
    process(s_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(s_in_buffer, konst_9359_wire_constant, tmp_var);
      BITSEL_u8_u1_9360_wire <= tmp_var; -- 
    end process;
    -- 
  end Block; -- data_path
  -- 
end Inv_Sbox_4_Volatile_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library work;
use work.ahir_system_global_package.all;
entity MUL2_Volatile is -- 
  port ( -- 
    mul_in : in  std_logic_vector(7 downto 0);
    mul_out : out  std_logic_vector(7 downto 0)-- 
  );
  -- 
end entity MUL2_Volatile;
architecture MUL2_Volatile_arch of MUL2_Volatile is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector(8-1 downto 0);
  signal default_zero_sig: std_logic;
  -- input port buffer signals
  signal mul_in_buffer :  std_logic_vector(7 downto 0);
  -- output port buffer signals
  signal mul_out_buffer :  std_logic_vector(7 downto 0);
  -- volatile/operator module components. 
  -- 
begin --  
  -- input handling ------------------------------------------------
  mul_in_buffer <= mul_in;
  -- output handling  -------------------------------------------------------
  mul_out <= mul_out_buffer;
  -- the control path --------------------------------------------------
  default_zero_sig <= '0';
  -- volatile module, no control path
  -- the data path
  data_path: Block -- 
    signal BITSEL_u8_u1_9380_wire : std_logic_vector(0 downto 0);
    signal R_mod_const_9382_wire_constant : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_9383_wire : std_logic_vector(7 downto 0);
    signal inx2_9376 : std_logic_vector(7 downto 0);
    signal konst_9374_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9379_wire_constant : std_logic_vector(7 downto 0);
    signal xxMUL2xxmod_const : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    R_mod_const_9382_wire_constant <= "00011011";
    konst_9374_wire_constant <= "00000001";
    konst_9379_wire_constant <= "00000111";
    xxMUL2xxmod_const <= "00011011";
    -- flow-through select operator MUX_9385_inst
    mul_out_buffer <= XOR_u8_u8_9383_wire when (BITSEL_u8_u1_9380_wire(0) /=  '0') else inx2_9376;
    -- binary operator BITSEL_u8_u1_9380_inst
    process(mul_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(mul_in_buffer, konst_9379_wire_constant, tmp_var);
      BITSEL_u8_u1_9380_wire <= tmp_var; -- 
    end process;
    -- binary operator SHL_u8_u8_9375_inst
    process(mul_in_buffer) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntSHL_proc(mul_in_buffer, konst_9374_wire_constant, tmp_var);
      inx2_9376 <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_9383_inst
    process(inx2_9376) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(inx2_9376, R_mod_const_9382_wire_constant, tmp_var);
      XOR_u8_u8_9383_wire <= tmp_var; -- 
    end process;
    -- 
  end Block; -- data_path
  -- 
end MUL2_Volatile_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library work;
use work.ahir_system_global_package.all;
entity Out_wrap_daemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    e_out_buf_pipe_read_req : out  std_logic_vector(0 downto 0);
    e_out_buf_pipe_read_ack : in   std_logic_vector(0 downto 0);
    e_out_buf_pipe_read_data : in   std_logic_vector(127 downto 0);
    d_out_buf_pipe_read_req : out  std_logic_vector(0 downto 0);
    d_out_buf_pipe_read_ack : in   std_logic_vector(0 downto 0);
    d_out_buf_pipe_read_data : in   std_logic_vector(127 downto 0);
    out_wrap_cmd_pipe_read_req : out  std_logic_vector(0 downto 0);
    out_wrap_cmd_pipe_read_ack : in   std_logic_vector(0 downto 0);
    out_wrap_cmd_pipe_read_data : in   std_logic_vector(63 downto 0);
    out_wrap_data_pipe_read_req : out  std_logic_vector(0 downto 0);
    out_wrap_data_pipe_read_ack : in   std_logic_vector(0 downto 0);
    out_wrap_data_pipe_read_data : in   std_logic_vector(127 downto 0);
    status_out_pipe_read_req : out  std_logic_vector(0 downto 0);
    status_out_pipe_read_ack : in   std_logic_vector(0 downto 0);
    status_out_pipe_read_data : in   std_logic_vector(63 downto 0);
    w_out_buf_pipe_write_req : out  std_logic_vector(0 downto 0);
    w_out_buf_pipe_write_ack : in   std_logic_vector(0 downto 0);
    w_out_buf_pipe_write_data : out  std_logic_vector(127 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity Out_wrap_daemon;
architecture Out_wrap_daemon_arch of Out_wrap_daemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal Out_wrap_daemon_CP_855_start: Boolean;
  signal Out_wrap_daemon_CP_855_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal RPIPE_e_out_buf_9459_inst_req_0 : boolean;
  signal WPIPE_w_out_buf_9458_inst_ack_0 : boolean;
  signal RPIPE_e_out_buf_9459_inst_ack_0 : boolean;
  signal OR_u15_u15_9446_inst_req_1 : boolean;
  signal WPIPE_w_out_buf_9458_inst_req_0 : boolean;
  signal RPIPE_out_wrap_data_9488_inst_req_1 : boolean;
  signal OR_u15_u15_9446_inst_ack_0 : boolean;
  signal RPIPE_d_out_buf_9463_inst_ack_0 : boolean;
  signal if_stmt_9471_branch_ack_0 : boolean;
  signal if_stmt_9454_branch_ack_1 : boolean;
  signal RPIPE_out_wrap_data_9488_inst_req_0 : boolean;
  signal WPIPE_w_out_buf_9462_inst_req_1 : boolean;
  signal if_stmt_9454_branch_ack_0 : boolean;
  signal WPIPE_w_out_buf_9462_inst_ack_1 : boolean;
  signal WPIPE_w_out_buf_9462_inst_req_0 : boolean;
  signal if_stmt_9477_branch_ack_1 : boolean;
  signal WPIPE_w_out_buf_9462_inst_ack_0 : boolean;
  signal OR_u15_u15_9446_inst_ack_1 : boolean;
  signal RPIPE_out_wrap_data_9488_inst_ack_1 : boolean;
  signal RPIPE_d_out_buf_9463_inst_req_0 : boolean;
  signal RPIPE_out_wrap_data_9488_inst_ack_0 : boolean;
  signal if_stmt_9477_branch_ack_0 : boolean;
  signal OR_u15_u15_9446_inst_req_0 : boolean;
  signal if_stmt_9477_branch_req_0 : boolean;
  signal RPIPE_e_out_buf_9459_inst_ack_1 : boolean;
  signal if_stmt_9454_branch_req_0 : boolean;
  signal RPIPE_out_wrap_cmd_9403_inst_req_0 : boolean;
  signal RPIPE_out_wrap_cmd_9403_inst_ack_0 : boolean;
  signal RPIPE_out_wrap_cmd_9403_inst_req_1 : boolean;
  signal RPIPE_out_wrap_cmd_9403_inst_ack_1 : boolean;
  signal if_stmt_9471_branch_ack_1 : boolean;
  signal RPIPE_status_out_9406_inst_req_0 : boolean;
  signal RPIPE_status_out_9406_inst_ack_0 : boolean;
  signal RPIPE_status_out_9406_inst_req_1 : boolean;
  signal RPIPE_status_out_9406_inst_ack_1 : boolean;
  signal if_stmt_9471_branch_req_0 : boolean;
  signal CONCAT_u64_u128_9411_inst_req_0 : boolean;
  signal CONCAT_u64_u128_9411_inst_ack_0 : boolean;
  signal CONCAT_u64_u128_9411_inst_req_1 : boolean;
  signal CONCAT_u64_u128_9411_inst_ack_1 : boolean;
  signal WPIPE_w_out_buf_9487_inst_req_0 : boolean;
  signal WPIPE_w_out_buf_9487_inst_ack_0 : boolean;
  signal WPIPE_w_out_buf_9408_inst_req_0 : boolean;
  signal WPIPE_w_out_buf_9408_inst_ack_0 : boolean;
  signal WPIPE_w_out_buf_9408_inst_req_1 : boolean;
  signal WPIPE_w_out_buf_9408_inst_ack_1 : boolean;
  signal WPIPE_w_out_buf_9458_inst_ack_1 : boolean;
  signal WPIPE_w_out_buf_9458_inst_req_1 : boolean;
  signal RPIPE_e_out_buf_9459_inst_req_1 : boolean;
  signal RPIPE_d_out_buf_9463_inst_ack_1 : boolean;
  signal RPIPE_d_out_buf_9463_inst_req_1 : boolean;
  signal WPIPE_w_out_buf_9487_inst_req_1 : boolean;
  signal WPIPE_w_out_buf_9487_inst_ack_1 : boolean;
  signal if_stmt_9495_branch_req_0 : boolean;
  signal if_stmt_9495_branch_ack_1 : boolean;
  signal if_stmt_9495_branch_ack_0 : boolean;
  signal n_count_var_9470_9484_buf_req_0 : boolean;
  signal n_count_var_9470_9484_buf_ack_0 : boolean;
  signal n_count_var_9470_9484_buf_req_1 : boolean;
  signal n_count_var_9470_9484_buf_ack_1 : boolean;
  signal phi_stmt_9482_req_0 : boolean;
  signal n_count_var2_9494_9485_buf_req_0 : boolean;
  signal n_count_var2_9494_9485_buf_ack_0 : boolean;
  signal n_count_var2_9494_9485_buf_req_1 : boolean;
  signal n_count_var2_9494_9485_buf_ack_1 : boolean;
  signal phi_stmt_9482_req_1 : boolean;
  signal phi_stmt_9482_ack_0 : boolean;
  signal phi_stmt_9449_req_0 : boolean;
  signal n_count_var_9470_9452_buf_req_0 : boolean;
  signal n_count_var_9470_9452_buf_ack_0 : boolean;
  signal n_count_var_9470_9452_buf_req_1 : boolean;
  signal n_count_var_9470_9452_buf_ack_1 : boolean;
  signal phi_stmt_9449_req_1 : boolean;
  signal phi_stmt_9449_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "Out_wrap_daemon_input_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      bypass_flag => true,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  Out_wrap_daemon_CP_855_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "Out_wrap_daemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= Out_wrap_daemon_CP_855_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= Out_wrap_daemon_CP_855_start & tag_ilock_write_ack_symbol;
    gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= Out_wrap_daemon_CP_855_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  Out_wrap_daemon_CP_855: Block -- control-path 
    signal Out_wrap_daemon_CP_855_elements: BooleanArray(103 downto 0);
    -- 
  begin -- 
    Out_wrap_daemon_CP_855_elements(0) <= Out_wrap_daemon_CP_855_start;
    Out_wrap_daemon_CP_855_symbol <= Out_wrap_daemon_CP_855_elements(103);
    -- CP-element group 0:  transition  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (2) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_9401/$entry
      -- 
    -- CP-element group 1:  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	9 
    -- CP-element group 1:  members (2) 
      -- CP-element group 1: 	 branch_block_stmt_9401/branch_block_stmt_9401__entry__
      -- CP-element group 1: 	 branch_block_stmt_9401/assign_stmt_9404__entry__
      -- 
    Out_wrap_daemon_CP_855_elements(1) <= Out_wrap_daemon_CP_855_elements(0);
    -- CP-element group 2:  place  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	11 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	12 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_9401/assign_stmt_9404__exit__
      -- CP-element group 2: 	 branch_block_stmt_9401/assign_stmt_9407__entry__
      -- 
    Out_wrap_daemon_CP_855_elements(2) <= Out_wrap_daemon_CP_855_elements(11);
    -- CP-element group 3:  place  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	14 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	15 
    -- CP-element group 3:  members (2) 
      -- CP-element group 3: 	 branch_block_stmt_9401/assign_stmt_9407__exit__
      -- CP-element group 3: 	 branch_block_stmt_9401/assign_stmt_9412__entry__
      -- 
    Out_wrap_daemon_CP_855_elements(3) <= Out_wrap_daemon_CP_855_elements(14);
    -- CP-element group 4:  place  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	19 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	20 
    -- CP-element group 4:  members (2) 
      -- CP-element group 4: 	 branch_block_stmt_9401/assign_stmt_9412__exit__
      -- CP-element group 4: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447__entry__
      -- 
    Out_wrap_daemon_CP_855_elements(4) <= Out_wrap_daemon_CP_855_elements(19);
    -- CP-element group 5:  branch  place  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	23 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	94 
    -- CP-element group 5: 	95 
    -- CP-element group 5:  members (2) 
      -- CP-element group 5: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447__exit__
      -- CP-element group 5: 	 branch_block_stmt_9401/merge_stmt_9448__entry__
      -- 
    Out_wrap_daemon_CP_855_elements(5) <= Out_wrap_daemon_CP_855_elements(23);
    -- CP-element group 6:  merge  branch  place  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	102 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	24 
    -- CP-element group 6: 	25 
    -- CP-element group 6:  members (2) 
      -- CP-element group 6: 	 branch_block_stmt_9401/merge_stmt_9448__exit__
      -- CP-element group 6: 	 branch_block_stmt_9401/if_stmt_9454__entry__
      -- 
    Out_wrap_daemon_CP_855_elements(6) <= Out_wrap_daemon_CP_855_elements(102);
    -- CP-element group 7:  merge  place  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	32 
    -- CP-element group 7: 	39 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	45 
    -- CP-element group 7:  members (2) 
      -- CP-element group 7: 	 branch_block_stmt_9401/if_stmt_9454__exit__
      -- CP-element group 7: 	 branch_block_stmt_9401/assign_stmt_9470__entry__
      -- 
    Out_wrap_daemon_CP_855_elements(7) <= OrReduce(Out_wrap_daemon_CP_855_elements(32) & Out_wrap_daemon_CP_855_elements(39));
    -- CP-element group 8:  branch  place  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	45 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	46 
    -- CP-element group 8: 	47 
    -- CP-element group 8:  members (2) 
      -- CP-element group 8: 	 branch_block_stmt_9401/assign_stmt_9470__exit__
      -- CP-element group 8: 	 branch_block_stmt_9401/if_stmt_9471__entry__
      -- 
    Out_wrap_daemon_CP_855_elements(8) <= Out_wrap_daemon_CP_855_elements(45);
    -- CP-element group 9:  transition  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	1 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (4) 
      -- CP-element group 9: 	 branch_block_stmt_9401/assign_stmt_9404/$entry
      -- CP-element group 9: 	 branch_block_stmt_9401/assign_stmt_9404/RPIPE_out_wrap_cmd_9403_sample_start_
      -- CP-element group 9: 	 branch_block_stmt_9401/assign_stmt_9404/RPIPE_out_wrap_cmd_9403_Sample/$entry
      -- CP-element group 9: 	 branch_block_stmt_9401/assign_stmt_9404/RPIPE_out_wrap_cmd_9403_Sample/rr
      -- 
    rr_889_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_889_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => Out_wrap_daemon_CP_855_elements(9), ack => RPIPE_out_wrap_cmd_9403_inst_req_0); -- 
    Out_wrap_daemon_CP_855_elements(9) <= Out_wrap_daemon_CP_855_elements(1);
    -- CP-element group 10:  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (6) 
      -- CP-element group 10: 	 branch_block_stmt_9401/assign_stmt_9404/RPIPE_out_wrap_cmd_9403_sample_completed_
      -- CP-element group 10: 	 branch_block_stmt_9401/assign_stmt_9404/RPIPE_out_wrap_cmd_9403_update_start_
      -- CP-element group 10: 	 branch_block_stmt_9401/assign_stmt_9404/RPIPE_out_wrap_cmd_9403_Sample/$exit
      -- CP-element group 10: 	 branch_block_stmt_9401/assign_stmt_9404/RPIPE_out_wrap_cmd_9403_Sample/ra
      -- CP-element group 10: 	 branch_block_stmt_9401/assign_stmt_9404/RPIPE_out_wrap_cmd_9403_Update/$entry
      -- CP-element group 10: 	 branch_block_stmt_9401/assign_stmt_9404/RPIPE_out_wrap_cmd_9403_Update/cr
      -- 
    ra_890_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_out_wrap_cmd_9403_inst_ack_0, ack => Out_wrap_daemon_CP_855_elements(10)); -- 
    cr_894_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_894_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => Out_wrap_daemon_CP_855_elements(10), ack => RPIPE_out_wrap_cmd_9403_inst_req_1); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	2 
    -- CP-element group 11:  members (4) 
      -- CP-element group 11: 	 branch_block_stmt_9401/assign_stmt_9404/$exit
      -- CP-element group 11: 	 branch_block_stmt_9401/assign_stmt_9404/RPIPE_out_wrap_cmd_9403_update_completed_
      -- CP-element group 11: 	 branch_block_stmt_9401/assign_stmt_9404/RPIPE_out_wrap_cmd_9403_Update/$exit
      -- CP-element group 11: 	 branch_block_stmt_9401/assign_stmt_9404/RPIPE_out_wrap_cmd_9403_Update/ca
      -- 
    ca_895_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_out_wrap_cmd_9403_inst_ack_1, ack => Out_wrap_daemon_CP_855_elements(11)); -- 
    -- CP-element group 12:  transition  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	2 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (4) 
      -- CP-element group 12: 	 branch_block_stmt_9401/assign_stmt_9407/$entry
      -- CP-element group 12: 	 branch_block_stmt_9401/assign_stmt_9407/RPIPE_status_out_9406_sample_start_
      -- CP-element group 12: 	 branch_block_stmt_9401/assign_stmt_9407/RPIPE_status_out_9406_Sample/$entry
      -- CP-element group 12: 	 branch_block_stmt_9401/assign_stmt_9407/RPIPE_status_out_9406_Sample/rr
      -- 
    rr_906_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_906_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => Out_wrap_daemon_CP_855_elements(12), ack => RPIPE_status_out_9406_inst_req_0); -- 
    Out_wrap_daemon_CP_855_elements(12) <= Out_wrap_daemon_CP_855_elements(2);
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_9401/assign_stmt_9407/RPIPE_status_out_9406_sample_completed_
      -- CP-element group 13: 	 branch_block_stmt_9401/assign_stmt_9407/RPIPE_status_out_9406_update_start_
      -- CP-element group 13: 	 branch_block_stmt_9401/assign_stmt_9407/RPIPE_status_out_9406_Sample/$exit
      -- CP-element group 13: 	 branch_block_stmt_9401/assign_stmt_9407/RPIPE_status_out_9406_Sample/ra
      -- CP-element group 13: 	 branch_block_stmt_9401/assign_stmt_9407/RPIPE_status_out_9406_Update/$entry
      -- CP-element group 13: 	 branch_block_stmt_9401/assign_stmt_9407/RPIPE_status_out_9406_Update/cr
      -- 
    ra_907_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_status_out_9406_inst_ack_0, ack => Out_wrap_daemon_CP_855_elements(13)); -- 
    cr_911_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_911_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => Out_wrap_daemon_CP_855_elements(13), ack => RPIPE_status_out_9406_inst_req_1); -- 
    -- CP-element group 14:  transition  input  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	3 
    -- CP-element group 14:  members (4) 
      -- CP-element group 14: 	 branch_block_stmt_9401/assign_stmt_9407/$exit
      -- CP-element group 14: 	 branch_block_stmt_9401/assign_stmt_9407/RPIPE_status_out_9406_update_completed_
      -- CP-element group 14: 	 branch_block_stmt_9401/assign_stmt_9407/RPIPE_status_out_9406_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_9401/assign_stmt_9407/RPIPE_status_out_9406_Update/ca
      -- 
    ca_912_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_status_out_9406_inst_ack_1, ack => Out_wrap_daemon_CP_855_elements(14)); -- 
    -- CP-element group 15:  join  fork  transition  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	3 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15: 	17 
    -- CP-element group 15:  members (15) 
      -- CP-element group 15: 	 branch_block_stmt_9401/assign_stmt_9412/$entry
      -- CP-element group 15: 	 branch_block_stmt_9401/assign_stmt_9412/CONCAT_u64_u128_9411_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_9401/assign_stmt_9412/CONCAT_u64_u128_9411_update_start_
      -- CP-element group 15: 	 branch_block_stmt_9401/assign_stmt_9412/R_head_out_9409_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_9401/assign_stmt_9412/R_head_out_9409_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_9401/assign_stmt_9412/R_head_out_9409_update_start_
      -- CP-element group 15: 	 branch_block_stmt_9401/assign_stmt_9412/R_head_out_9409_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_9401/assign_stmt_9412/R_st_out_9410_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_9401/assign_stmt_9412/R_st_out_9410_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_9401/assign_stmt_9412/R_st_out_9410_update_start_
      -- CP-element group 15: 	 branch_block_stmt_9401/assign_stmt_9412/R_st_out_9410_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_9401/assign_stmt_9412/CONCAT_u64_u128_9411_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_9401/assign_stmt_9412/CONCAT_u64_u128_9411_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_9401/assign_stmt_9412/CONCAT_u64_u128_9411_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_9401/assign_stmt_9412/CONCAT_u64_u128_9411_Update/cr
      -- 
    cr_936_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_936_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => Out_wrap_daemon_CP_855_elements(15), ack => CONCAT_u64_u128_9411_inst_req_1); -- 
    rr_931_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_931_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => Out_wrap_daemon_CP_855_elements(15), ack => CONCAT_u64_u128_9411_inst_req_0); -- 
    Out_wrap_daemon_CP_855_elements(15) <= Out_wrap_daemon_CP_855_elements(3);
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_9401/assign_stmt_9412/CONCAT_u64_u128_9411_sample_completed_
      -- CP-element group 16: 	 branch_block_stmt_9401/assign_stmt_9412/CONCAT_u64_u128_9411_Sample/$exit
      -- CP-element group 16: 	 branch_block_stmt_9401/assign_stmt_9412/CONCAT_u64_u128_9411_Sample/ra
      -- 
    ra_932_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u64_u128_9411_inst_ack_0, ack => Out_wrap_daemon_CP_855_elements(16)); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	15 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_9401/assign_stmt_9412/CONCAT_u64_u128_9411_update_completed_
      -- CP-element group 17: 	 branch_block_stmt_9401/assign_stmt_9412/CONCAT_u64_u128_9411_Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_9401/assign_stmt_9412/CONCAT_u64_u128_9411_Update/ca
      -- CP-element group 17: 	 branch_block_stmt_9401/assign_stmt_9412/WPIPE_w_out_buf_9408_sample_start_
      -- CP-element group 17: 	 branch_block_stmt_9401/assign_stmt_9412/WPIPE_w_out_buf_9408_Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_9401/assign_stmt_9412/WPIPE_w_out_buf_9408_Sample/req
      -- 
    ca_937_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u64_u128_9411_inst_ack_1, ack => Out_wrap_daemon_CP_855_elements(17)); -- 
    req_945_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_945_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => Out_wrap_daemon_CP_855_elements(17), ack => WPIPE_w_out_buf_9408_inst_req_0); -- 
    -- CP-element group 18:  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (6) 
      -- CP-element group 18: 	 branch_block_stmt_9401/assign_stmt_9412/WPIPE_w_out_buf_9408_sample_completed_
      -- CP-element group 18: 	 branch_block_stmt_9401/assign_stmt_9412/WPIPE_w_out_buf_9408_update_start_
      -- CP-element group 18: 	 branch_block_stmt_9401/assign_stmt_9412/WPIPE_w_out_buf_9408_Sample/$exit
      -- CP-element group 18: 	 branch_block_stmt_9401/assign_stmt_9412/WPIPE_w_out_buf_9408_Sample/ack
      -- CP-element group 18: 	 branch_block_stmt_9401/assign_stmt_9412/WPIPE_w_out_buf_9408_Update/$entry
      -- CP-element group 18: 	 branch_block_stmt_9401/assign_stmt_9412/WPIPE_w_out_buf_9408_Update/req
      -- 
    ack_946_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_w_out_buf_9408_inst_ack_0, ack => Out_wrap_daemon_CP_855_elements(18)); -- 
    req_950_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_950_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => Out_wrap_daemon_CP_855_elements(18), ack => WPIPE_w_out_buf_9408_inst_req_1); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	4 
    -- CP-element group 19:  members (4) 
      -- CP-element group 19: 	 branch_block_stmt_9401/assign_stmt_9412/$exit
      -- CP-element group 19: 	 branch_block_stmt_9401/assign_stmt_9412/WPIPE_w_out_buf_9408_update_completed_
      -- CP-element group 19: 	 branch_block_stmt_9401/assign_stmt_9412/WPIPE_w_out_buf_9408_Update/$exit
      -- CP-element group 19: 	 branch_block_stmt_9401/assign_stmt_9412/WPIPE_w_out_buf_9408_Update/ack
      -- 
    ack_951_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_w_out_buf_9408_inst_ack_1, ack => Out_wrap_daemon_CP_855_elements(19)); -- 
    -- CP-element group 20:  join  fork  transition  output  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	4 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	21 
    -- CP-element group 20: 	22 
    -- CP-element group 20: 	23 
    -- CP-element group 20:  members (147) 
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/R_count_9435_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/UGE_u15_u1_9442_Sample/ra
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/R_count_9435_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/R_count_9441_sample_start_
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/ULT_u15_u1_9436_Update/cr
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/ULT_u15_u1_9436_Update/ca
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/ULT_u15_u1_9436_Sample/$entry
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/UGE_u15_u1_9442_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/R_count_9435_update_start_
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/UGE_u15_u1_9442_Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/UGE_u15_u1_9442_Update/$entry
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/OR_u15_u15_9446_Update/cr
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/UGE_u15_u1_9442_update_start_
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/UGE_u15_u1_9442_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/ULT_u15_u1_9436_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/UGE_u15_u1_9442_sample_start_
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/OR_u15_u15_9446_Update/$entry
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/MUX_9445_complete/$exit
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/R_count_9443_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/MUX_9445_complete/req
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/MUX_9439_start/$entry
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/MUX_9439_start/$exit
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/MUX_9439_start/req
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/R_count_9443_update_start_
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/R_count_9443_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/MUX_9445_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/MUX_9445_start/$entry
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/MUX_9439_start/ack
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/R_count_9441_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/MUX_9445_complete/ack
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/MUX_9439_complete/$entry
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/ULT_u15_u1_9436_Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/MUX_9445_start/$exit
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/MUX_9445_start/req
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/UGE_u15_u1_9442_Sample/rr
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/MUX_9439_complete/$exit
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/UGE_u15_u1_9442_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/R_count_9441_update_start_
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/UGE_u15_u1_9442_Update/cr
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/MUX_9439_complete/req
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/MUX_9439_complete/ack
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/MUX_9445_sample_start_
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/MUX_9445_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/MUX_9445_update_start_
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/MUX_9445_start/ack
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/R_count_9441_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/MUX_9445_complete/$entry
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/UGE_u15_u1_9442_Sample/$entry
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/UGE_u15_u1_9442_Update/ca
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/OR_u15_u15_9446_Sample/rr
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/ULT_u15_u1_9436_Update/$entry
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/ULT_u15_u1_9436_Sample/ra
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/ULT_u15_u1_9436_Sample/rr
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/R_count_9435_sample_start_
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/ULT_u15_u1_9436_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/ULT_u15_u1_9436_update_start_
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/$entry
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/slice_9415_sample_start_
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/slice_9415_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/slice_9415_update_start_
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/slice_9415_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/R_head_out_9414_sample_start_
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/R_head_out_9414_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/R_head_out_9414_update_start_
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/R_head_out_9414_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/slice_9415_Sample/$entry
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/slice_9415_Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/slice_9415_Sample/rr
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/slice_9415_Sample/ra
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/OR_u15_u15_9446_Sample/$entry
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/slice_9415_Update/$entry
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/slice_9415_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/slice_9415_Update/cr
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/slice_9415_Update/ca
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/slice_9419_sample_start_
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/slice_9419_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/slice_9419_update_start_
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/slice_9419_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/R_head_out_9418_sample_start_
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/R_head_out_9418_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/R_head_out_9418_update_start_
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/R_head_out_9418_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/slice_9419_Sample/$entry
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/slice_9419_Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/slice_9419_Sample/rr
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/slice_9419_Sample/ra
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/slice_9419_Update/$entry
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/slice_9419_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/slice_9419_Update/cr
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/slice_9419_Update/ca
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/slice_9423_sample_start_
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/slice_9423_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/slice_9423_update_start_
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/slice_9423_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/R_head_out_9422_sample_start_
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/R_head_out_9422_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/R_head_out_9422_update_start_
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/R_head_out_9422_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/slice_9423_Sample/$entry
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/slice_9423_Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/slice_9423_Sample/rr
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/slice_9423_Sample/ra
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/slice_9423_Update/$entry
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/slice_9423_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/slice_9423_Update/cr
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/slice_9423_Update/ca
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/slice_9427_sample_start_
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/slice_9427_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/slice_9427_update_start_
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/slice_9427_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/R_head_out_9426_sample_start_
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/R_head_out_9426_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/R_head_out_9426_update_start_
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/R_head_out_9426_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/slice_9427_Sample/$entry
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/slice_9427_Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/slice_9427_Sample/rr
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/slice_9427_Sample/ra
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/slice_9427_Update/$entry
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/slice_9427_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/R_count_9443_sample_start_
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/slice_9427_Update/cr
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/slice_9427_Update/ca
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/slice_9431_sample_start_
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/slice_9431_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/slice_9431_update_start_
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/slice_9431_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/R_head_out_9430_sample_start_
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/R_head_out_9430_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/R_head_out_9430_update_start_
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/R_head_out_9430_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/slice_9431_Sample/$entry
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/slice_9431_Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/slice_9431_Sample/rr
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/slice_9431_Sample/ra
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/slice_9431_Update/$entry
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/slice_9431_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/slice_9431_Update/cr
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/slice_9431_Update/ca
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/OR_u15_u15_9446_sample_start_
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/OR_u15_u15_9446_update_start_
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/MUX_9439_sample_start_
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/MUX_9439_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/MUX_9439_update_start_
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/MUX_9439_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/ULT_u15_u1_9436_sample_start_
      -- CP-element group 20: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/ULT_u15_u1_9436_sample_completed_
      -- 
    rr_1120_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1120_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => Out_wrap_daemon_CP_855_elements(20), ack => OR_u15_u15_9446_inst_req_0); -- 
    cr_1125_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1125_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => Out_wrap_daemon_CP_855_elements(20), ack => OR_u15_u15_9446_inst_req_1); -- 
    Out_wrap_daemon_CP_855_elements(20) <= Out_wrap_daemon_CP_855_elements(4);
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	20 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/OR_u15_u15_9446_Sample/ra
      -- CP-element group 21: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/OR_u15_u15_9446_Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/OR_u15_u15_9446_sample_completed_
      -- 
    ra_1121_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => OR_u15_u15_9446_inst_ack_0, ack => Out_wrap_daemon_CP_855_elements(21)); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	20 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	23 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/OR_u15_u15_9446_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/OR_u15_u15_9446_Update/ca
      -- CP-element group 22: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/OR_u15_u15_9446_update_completed_
      -- 
    ca_1126_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => OR_u15_u15_9446_inst_ack_1, ack => Out_wrap_daemon_CP_855_elements(22)); -- 
    -- CP-element group 23:  join  transition  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	20 
    -- CP-element group 23: 	22 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	5 
    -- CP-element group 23:  members (1) 
      -- CP-element group 23: 	 branch_block_stmt_9401/assign_stmt_9416_to_assign_stmt_9447/$exit
      -- 
    Out_wrap_daemon_cp_element_group_23: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "Out_wrap_daemon_cp_element_group_23"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= Out_wrap_daemon_CP_855_elements(20) & Out_wrap_daemon_CP_855_elements(22);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => Out_wrap_daemon_CP_855_elements(23), clk => clk, reset => reset); --
    end block;
    -- CP-element group 24:  transition  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	6 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (1) 
      -- CP-element group 24: 	 branch_block_stmt_9401/if_stmt_9454_dead_link/$entry
      -- 
    Out_wrap_daemon_CP_855_elements(24) <= Out_wrap_daemon_CP_855_elements(6);
    -- CP-element group 25:  transition  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	6 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25:  members (17) 
      -- CP-element group 25: 	 branch_block_stmt_9401/if_stmt_9454_eval_test/branch_req
      -- CP-element group 25: 	 branch_block_stmt_9401/if_stmt_9454_eval_test/EQ_u1_u1_9457/SplitProtocol/Update/ca
      -- CP-element group 25: 	 branch_block_stmt_9401/if_stmt_9454_eval_test/EQ_u1_u1_9457/SplitProtocol/Update/cr
      -- CP-element group 25: 	 branch_block_stmt_9401/if_stmt_9454_eval_test/EQ_u1_u1_9457/SplitProtocol/Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_9401/if_stmt_9454_eval_test/EQ_u1_u1_9457/SplitProtocol/Update/$entry
      -- CP-element group 25: 	 branch_block_stmt_9401/if_stmt_9454_eval_test/EQ_u1_u1_9457/SplitProtocol/Sample/ra
      -- CP-element group 25: 	 branch_block_stmt_9401/if_stmt_9454_eval_test/EQ_u1_u1_9457/SplitProtocol/Sample/rr
      -- CP-element group 25: 	 branch_block_stmt_9401/if_stmt_9454_eval_test/EQ_u1_u1_9457/SplitProtocol/Sample/$exit
      -- CP-element group 25: 	 branch_block_stmt_9401/if_stmt_9454_eval_test/EQ_u1_u1_9457/SplitProtocol/Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_9401/if_stmt_9454_eval_test/EQ_u1_u1_9457/SplitProtocol/$exit
      -- CP-element group 25: 	 branch_block_stmt_9401/if_stmt_9454_eval_test/EQ_u1_u1_9457/SplitProtocol/$entry
      -- CP-element group 25: 	 branch_block_stmt_9401/if_stmt_9454_eval_test/EQ_u1_u1_9457/EQ_u1_u1_9457_inputs/$exit
      -- CP-element group 25: 	 branch_block_stmt_9401/if_stmt_9454_eval_test/EQ_u1_u1_9457/EQ_u1_u1_9457_inputs/$entry
      -- CP-element group 25: 	 branch_block_stmt_9401/if_stmt_9454_eval_test/EQ_u1_u1_9457/$exit
      -- CP-element group 25: 	 branch_block_stmt_9401/if_stmt_9454_eval_test/EQ_u1_u1_9457/$entry
      -- CP-element group 25: 	 branch_block_stmt_9401/if_stmt_9454_eval_test/$exit
      -- CP-element group 25: 	 branch_block_stmt_9401/if_stmt_9454_eval_test/$entry
      -- 
    branch_req_1153_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1153_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => Out_wrap_daemon_CP_855_elements(25), ack => if_stmt_9454_branch_req_0); -- 
    Out_wrap_daemon_CP_855_elements(25) <= Out_wrap_daemon_CP_855_elements(6);
    -- CP-element group 26:  branch  place  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	25 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	27 
    -- CP-element group 26: 	29 
    -- CP-element group 26:  members (1) 
      -- CP-element group 26: 	 branch_block_stmt_9401/EQ_u1_u1_9457_place
      -- 
    Out_wrap_daemon_CP_855_elements(26) <= Out_wrap_daemon_CP_855_elements(25);
    -- CP-element group 27:  transition  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	26 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	28 
    -- CP-element group 27:  members (1) 
      -- CP-element group 27: 	 branch_block_stmt_9401/if_stmt_9454_if_link/$entry
      -- 
    Out_wrap_daemon_CP_855_elements(27) <= Out_wrap_daemon_CP_855_elements(26);
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	27 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	31 
    -- CP-element group 28:  members (2) 
      -- CP-element group 28: 	 branch_block_stmt_9401/if_stmt_9454_if_link/$exit
      -- CP-element group 28: 	 branch_block_stmt_9401/if_stmt_9454_if_link/if_choice_transition
      -- 
    if_choice_transition_1158_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_9454_branch_ack_1, ack => Out_wrap_daemon_CP_855_elements(28)); -- 
    -- CP-element group 29:  transition  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	26 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (1) 
      -- CP-element group 29: 	 branch_block_stmt_9401/if_stmt_9454_else_link/$entry
      -- 
    Out_wrap_daemon_CP_855_elements(29) <= Out_wrap_daemon_CP_855_elements(26);
    -- CP-element group 30:  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	38 
    -- CP-element group 30:  members (2) 
      -- CP-element group 30: 	 branch_block_stmt_9401/if_stmt_9454_else_link/$exit
      -- CP-element group 30: 	 branch_block_stmt_9401/if_stmt_9454_else_link/else_choice_transition
      -- 
    else_choice_transition_1162_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_9454_branch_ack_0, ack => Out_wrap_daemon_CP_855_elements(30)); -- 
    -- CP-element group 31:  place  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	28 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	33 
    -- CP-element group 31:  members (1) 
      -- CP-element group 31: 	 branch_block_stmt_9401/assign_stmt_9460__entry__
      -- 
    Out_wrap_daemon_CP_855_elements(31) <= Out_wrap_daemon_CP_855_elements(28);
    -- CP-element group 32:  place  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	37 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	7 
    -- CP-element group 32:  members (1) 
      -- CP-element group 32: 	 branch_block_stmt_9401/assign_stmt_9460__exit__
      -- 
    Out_wrap_daemon_CP_855_elements(32) <= Out_wrap_daemon_CP_855_elements(37);
    -- CP-element group 33:  transition  output  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	31 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (4) 
      -- CP-element group 33: 	 branch_block_stmt_9401/assign_stmt_9460/RPIPE_e_out_buf_9459_Sample/rr
      -- CP-element group 33: 	 branch_block_stmt_9401/assign_stmt_9460/$entry
      -- CP-element group 33: 	 branch_block_stmt_9401/assign_stmt_9460/RPIPE_e_out_buf_9459_sample_start_
      -- CP-element group 33: 	 branch_block_stmt_9401/assign_stmt_9460/RPIPE_e_out_buf_9459_Sample/$entry
      -- 
    rr_1175_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1175_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => Out_wrap_daemon_CP_855_elements(33), ack => RPIPE_e_out_buf_9459_inst_req_0); -- 
    Out_wrap_daemon_CP_855_elements(33) <= Out_wrap_daemon_CP_855_elements(31);
    -- CP-element group 34:  transition  input  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34:  members (6) 
      -- CP-element group 34: 	 branch_block_stmt_9401/assign_stmt_9460/RPIPE_e_out_buf_9459_Sample/$exit
      -- CP-element group 34: 	 branch_block_stmt_9401/assign_stmt_9460/RPIPE_e_out_buf_9459_Sample/ra
      -- CP-element group 34: 	 branch_block_stmt_9401/assign_stmt_9460/RPIPE_e_out_buf_9459_sample_completed_
      -- CP-element group 34: 	 branch_block_stmt_9401/assign_stmt_9460/RPIPE_e_out_buf_9459_update_start_
      -- CP-element group 34: 	 branch_block_stmt_9401/assign_stmt_9460/RPIPE_e_out_buf_9459_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_9401/assign_stmt_9460/RPIPE_e_out_buf_9459_Update/$entry
      -- 
    ra_1176_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_e_out_buf_9459_inst_ack_0, ack => Out_wrap_daemon_CP_855_elements(34)); -- 
    cr_1180_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1180_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => Out_wrap_daemon_CP_855_elements(34), ack => RPIPE_e_out_buf_9459_inst_req_1); -- 
    -- CP-element group 35:  transition  input  output  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	36 
    -- CP-element group 35:  members (6) 
      -- CP-element group 35: 	 branch_block_stmt_9401/assign_stmt_9460/WPIPE_w_out_buf_9458_Sample/req
      -- CP-element group 35: 	 branch_block_stmt_9401/assign_stmt_9460/WPIPE_w_out_buf_9458_Sample/$entry
      -- CP-element group 35: 	 branch_block_stmt_9401/assign_stmt_9460/RPIPE_e_out_buf_9459_update_completed_
      -- CP-element group 35: 	 branch_block_stmt_9401/assign_stmt_9460/WPIPE_w_out_buf_9458_sample_start_
      -- CP-element group 35: 	 branch_block_stmt_9401/assign_stmt_9460/RPIPE_e_out_buf_9459_Update/ca
      -- CP-element group 35: 	 branch_block_stmt_9401/assign_stmt_9460/RPIPE_e_out_buf_9459_Update/$exit
      -- 
    ca_1181_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_e_out_buf_9459_inst_ack_1, ack => Out_wrap_daemon_CP_855_elements(35)); -- 
    req_1189_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1189_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => Out_wrap_daemon_CP_855_elements(35), ack => WPIPE_w_out_buf_9458_inst_req_0); -- 
    -- CP-element group 36:  transition  input  output  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	35 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	37 
    -- CP-element group 36:  members (6) 
      -- CP-element group 36: 	 branch_block_stmt_9401/assign_stmt_9460/WPIPE_w_out_buf_9458_Update/$entry
      -- CP-element group 36: 	 branch_block_stmt_9401/assign_stmt_9460/WPIPE_w_out_buf_9458_update_start_
      -- CP-element group 36: 	 branch_block_stmt_9401/assign_stmt_9460/WPIPE_w_out_buf_9458_Sample/ack
      -- CP-element group 36: 	 branch_block_stmt_9401/assign_stmt_9460/WPIPE_w_out_buf_9458_sample_completed_
      -- CP-element group 36: 	 branch_block_stmt_9401/assign_stmt_9460/WPIPE_w_out_buf_9458_Sample/$exit
      -- CP-element group 36: 	 branch_block_stmt_9401/assign_stmt_9460/WPIPE_w_out_buf_9458_Update/req
      -- 
    ack_1190_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_w_out_buf_9458_inst_ack_0, ack => Out_wrap_daemon_CP_855_elements(36)); -- 
    req_1194_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1194_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => Out_wrap_daemon_CP_855_elements(36), ack => WPIPE_w_out_buf_9458_inst_req_1); -- 
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	36 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	32 
    -- CP-element group 37:  members (4) 
      -- CP-element group 37: 	 branch_block_stmt_9401/assign_stmt_9460/WPIPE_w_out_buf_9458_update_completed_
      -- CP-element group 37: 	 branch_block_stmt_9401/assign_stmt_9460/$exit
      -- CP-element group 37: 	 branch_block_stmt_9401/assign_stmt_9460/WPIPE_w_out_buf_9458_Update/ack
      -- CP-element group 37: 	 branch_block_stmt_9401/assign_stmt_9460/WPIPE_w_out_buf_9458_Update/$exit
      -- 
    ack_1195_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_w_out_buf_9458_inst_ack_1, ack => Out_wrap_daemon_CP_855_elements(37)); -- 
    -- CP-element group 38:  place  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	30 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	40 
    -- CP-element group 38:  members (1) 
      -- CP-element group 38: 	 branch_block_stmt_9401/assign_stmt_9464__entry__
      -- 
    Out_wrap_daemon_CP_855_elements(38) <= Out_wrap_daemon_CP_855_elements(30);
    -- CP-element group 39:  place  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	44 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	7 
    -- CP-element group 39:  members (1) 
      -- CP-element group 39: 	 branch_block_stmt_9401/assign_stmt_9464__exit__
      -- 
    Out_wrap_daemon_CP_855_elements(39) <= Out_wrap_daemon_CP_855_elements(44);
    -- CP-element group 40:  transition  output  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	38 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	41 
    -- CP-element group 40:  members (4) 
      -- CP-element group 40: 	 branch_block_stmt_9401/assign_stmt_9464/RPIPE_d_out_buf_9463_Sample/$entry
      -- CP-element group 40: 	 branch_block_stmt_9401/assign_stmt_9464/RPIPE_d_out_buf_9463_sample_start_
      -- CP-element group 40: 	 branch_block_stmt_9401/assign_stmt_9464/RPIPE_d_out_buf_9463_Sample/rr
      -- CP-element group 40: 	 branch_block_stmt_9401/assign_stmt_9464/$entry
      -- 
    rr_1208_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1208_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => Out_wrap_daemon_CP_855_elements(40), ack => RPIPE_d_out_buf_9463_inst_req_0); -- 
    Out_wrap_daemon_CP_855_elements(40) <= Out_wrap_daemon_CP_855_elements(38);
    -- CP-element group 41:  transition  input  output  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	40 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	42 
    -- CP-element group 41:  members (6) 
      -- CP-element group 41: 	 branch_block_stmt_9401/assign_stmt_9464/RPIPE_d_out_buf_9463_sample_completed_
      -- CP-element group 41: 	 branch_block_stmt_9401/assign_stmt_9464/RPIPE_d_out_buf_9463_Sample/ra
      -- CP-element group 41: 	 branch_block_stmt_9401/assign_stmt_9464/RPIPE_d_out_buf_9463_Sample/$exit
      -- CP-element group 41: 	 branch_block_stmt_9401/assign_stmt_9464/RPIPE_d_out_buf_9463_Update/$entry
      -- CP-element group 41: 	 branch_block_stmt_9401/assign_stmt_9464/RPIPE_d_out_buf_9463_update_start_
      -- CP-element group 41: 	 branch_block_stmt_9401/assign_stmt_9464/RPIPE_d_out_buf_9463_Update/cr
      -- 
    ra_1209_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_d_out_buf_9463_inst_ack_0, ack => Out_wrap_daemon_CP_855_elements(41)); -- 
    cr_1213_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1213_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => Out_wrap_daemon_CP_855_elements(41), ack => RPIPE_d_out_buf_9463_inst_req_1); -- 
    -- CP-element group 42:  transition  input  output  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	41 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (6) 
      -- CP-element group 42: 	 branch_block_stmt_9401/assign_stmt_9464/WPIPE_w_out_buf_9462_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_9401/assign_stmt_9464/WPIPE_w_out_buf_9462_Sample/req
      -- CP-element group 42: 	 branch_block_stmt_9401/assign_stmt_9464/RPIPE_d_out_buf_9463_Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_9401/assign_stmt_9464/RPIPE_d_out_buf_9463_update_completed_
      -- CP-element group 42: 	 branch_block_stmt_9401/assign_stmt_9464/WPIPE_w_out_buf_9462_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_9401/assign_stmt_9464/RPIPE_d_out_buf_9463_Update/ca
      -- 
    ca_1214_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_d_out_buf_9463_inst_ack_1, ack => Out_wrap_daemon_CP_855_elements(42)); -- 
    req_1222_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1222_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => Out_wrap_daemon_CP_855_elements(42), ack => WPIPE_w_out_buf_9462_inst_req_0); -- 
    -- CP-element group 43:  transition  input  output  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	44 
    -- CP-element group 43:  members (6) 
      -- CP-element group 43: 	 branch_block_stmt_9401/assign_stmt_9464/WPIPE_w_out_buf_9462_Sample/$exit
      -- CP-element group 43: 	 branch_block_stmt_9401/assign_stmt_9464/WPIPE_w_out_buf_9462_update_start_
      -- CP-element group 43: 	 branch_block_stmt_9401/assign_stmt_9464/WPIPE_w_out_buf_9462_Update/$entry
      -- CP-element group 43: 	 branch_block_stmt_9401/assign_stmt_9464/WPIPE_w_out_buf_9462_Update/req
      -- CP-element group 43: 	 branch_block_stmt_9401/assign_stmt_9464/WPIPE_w_out_buf_9462_Sample/ack
      -- CP-element group 43: 	 branch_block_stmt_9401/assign_stmt_9464/WPIPE_w_out_buf_9462_sample_completed_
      -- 
    ack_1223_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_w_out_buf_9462_inst_ack_0, ack => Out_wrap_daemon_CP_855_elements(43)); -- 
    req_1227_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1227_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => Out_wrap_daemon_CP_855_elements(43), ack => WPIPE_w_out_buf_9462_inst_req_1); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	43 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	39 
    -- CP-element group 44:  members (4) 
      -- CP-element group 44: 	 branch_block_stmt_9401/assign_stmt_9464/WPIPE_w_out_buf_9462_update_completed_
      -- CP-element group 44: 	 branch_block_stmt_9401/assign_stmt_9464/WPIPE_w_out_buf_9462_Update/$exit
      -- CP-element group 44: 	 branch_block_stmt_9401/assign_stmt_9464/WPIPE_w_out_buf_9462_Update/ack
      -- CP-element group 44: 	 branch_block_stmt_9401/assign_stmt_9464/$exit
      -- 
    ack_1228_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_w_out_buf_9462_inst_ack_1, ack => Out_wrap_daemon_CP_855_elements(44)); -- 
    -- CP-element group 45:  transition  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	7 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	8 
    -- CP-element group 45:  members (18) 
      -- CP-element group 45: 	 branch_block_stmt_9401/assign_stmt_9470/R_count_var_9467_update_completed_
      -- CP-element group 45: 	 branch_block_stmt_9401/assign_stmt_9470/ADD_u15_u15_9469_Sample/$entry
      -- CP-element group 45: 	 branch_block_stmt_9401/assign_stmt_9470/R_count_var_9467_sample_start_
      -- CP-element group 45: 	 branch_block_stmt_9401/assign_stmt_9470/R_count_var_9467_sample_completed_
      -- CP-element group 45: 	 branch_block_stmt_9401/assign_stmt_9470/ADD_u15_u15_9469_Sample/$exit
      -- CP-element group 45: 	 branch_block_stmt_9401/assign_stmt_9470/R_count_var_9467_update_start_
      -- CP-element group 45: 	 branch_block_stmt_9401/assign_stmt_9470/$entry
      -- CP-element group 45: 	 branch_block_stmt_9401/assign_stmt_9470/$exit
      -- CP-element group 45: 	 branch_block_stmt_9401/assign_stmt_9470/ADD_u15_u15_9469_update_completed_
      -- CP-element group 45: 	 branch_block_stmt_9401/assign_stmt_9470/ADD_u15_u15_9469_update_start_
      -- CP-element group 45: 	 branch_block_stmt_9401/assign_stmt_9470/ADD_u15_u15_9469_sample_start_
      -- CP-element group 45: 	 branch_block_stmt_9401/assign_stmt_9470/ADD_u15_u15_9469_Update/ca
      -- CP-element group 45: 	 branch_block_stmt_9401/assign_stmt_9470/ADD_u15_u15_9469_Update/cr
      -- CP-element group 45: 	 branch_block_stmt_9401/assign_stmt_9470/ADD_u15_u15_9469_Update/$exit
      -- CP-element group 45: 	 branch_block_stmt_9401/assign_stmt_9470/ADD_u15_u15_9469_Update/$entry
      -- CP-element group 45: 	 branch_block_stmt_9401/assign_stmt_9470/ADD_u15_u15_9469_Sample/ra
      -- CP-element group 45: 	 branch_block_stmt_9401/assign_stmt_9470/ADD_u15_u15_9469_Sample/rr
      -- CP-element group 45: 	 branch_block_stmt_9401/assign_stmt_9470/ADD_u15_u15_9469_sample_completed_
      -- 
    Out_wrap_daemon_CP_855_elements(45) <= Out_wrap_daemon_CP_855_elements(7);
    -- CP-element group 46:  transition  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	8 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (1) 
      -- CP-element group 46: 	 branch_block_stmt_9401/if_stmt_9471_dead_link/$entry
      -- 
    Out_wrap_daemon_CP_855_elements(46) <= Out_wrap_daemon_CP_855_elements(8);
    -- CP-element group 47:  transition  output  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	8 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	48 
    -- CP-element group 47:  members (17) 
      -- CP-element group 47: 	 branch_block_stmt_9401/if_stmt_9471_eval_test/$entry
      -- CP-element group 47: 	 branch_block_stmt_9401/if_stmt_9471_eval_test/$exit
      -- CP-element group 47: 	 branch_block_stmt_9401/if_stmt_9471_eval_test/branch_req
      -- CP-element group 47: 	 branch_block_stmt_9401/if_stmt_9471_eval_test/ULT_u15_u1_9474/SplitProtocol/Update/ca
      -- CP-element group 47: 	 branch_block_stmt_9401/if_stmt_9471_eval_test/ULT_u15_u1_9474/SplitProtocol/Update/cr
      -- CP-element group 47: 	 branch_block_stmt_9401/if_stmt_9471_eval_test/ULT_u15_u1_9474/SplitProtocol/Update/$exit
      -- CP-element group 47: 	 branch_block_stmt_9401/if_stmt_9471_eval_test/ULT_u15_u1_9474/SplitProtocol/Update/$entry
      -- CP-element group 47: 	 branch_block_stmt_9401/if_stmt_9471_eval_test/ULT_u15_u1_9474/SplitProtocol/Sample/ra
      -- CP-element group 47: 	 branch_block_stmt_9401/if_stmt_9471_eval_test/ULT_u15_u1_9474/SplitProtocol/Sample/rr
      -- CP-element group 47: 	 branch_block_stmt_9401/if_stmt_9471_eval_test/ULT_u15_u1_9474/SplitProtocol/Sample/$exit
      -- CP-element group 47: 	 branch_block_stmt_9401/if_stmt_9471_eval_test/ULT_u15_u1_9474/SplitProtocol/Sample/$entry
      -- CP-element group 47: 	 branch_block_stmt_9401/if_stmt_9471_eval_test/ULT_u15_u1_9474/SplitProtocol/$exit
      -- CP-element group 47: 	 branch_block_stmt_9401/if_stmt_9471_eval_test/ULT_u15_u1_9474/SplitProtocol/$entry
      -- CP-element group 47: 	 branch_block_stmt_9401/if_stmt_9471_eval_test/ULT_u15_u1_9474/ULT_u15_u1_9474_inputs/$exit
      -- CP-element group 47: 	 branch_block_stmt_9401/if_stmt_9471_eval_test/ULT_u15_u1_9474/ULT_u15_u1_9474_inputs/$entry
      -- CP-element group 47: 	 branch_block_stmt_9401/if_stmt_9471_eval_test/ULT_u15_u1_9474/$exit
      -- CP-element group 47: 	 branch_block_stmt_9401/if_stmt_9471_eval_test/ULT_u15_u1_9474/$entry
      -- 
    branch_req_1276_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1276_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => Out_wrap_daemon_CP_855_elements(47), ack => if_stmt_9471_branch_req_0); -- 
    Out_wrap_daemon_CP_855_elements(47) <= Out_wrap_daemon_CP_855_elements(8);
    -- CP-element group 48:  branch  place  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	47 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	49 
    -- CP-element group 48: 	51 
    -- CP-element group 48:  members (1) 
      -- CP-element group 48: 	 branch_block_stmt_9401/ULT_u15_u1_9474_place
      -- 
    Out_wrap_daemon_CP_855_elements(48) <= Out_wrap_daemon_CP_855_elements(47);
    -- CP-element group 49:  transition  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	48 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (1) 
      -- CP-element group 49: 	 branch_block_stmt_9401/if_stmt_9471_if_link/$entry
      -- 
    Out_wrap_daemon_CP_855_elements(49) <= Out_wrap_daemon_CP_855_elements(48);
    -- CP-element group 50:  transition  input  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	53 
    -- CP-element group 50:  members (2) 
      -- CP-element group 50: 	 branch_block_stmt_9401/if_stmt_9471_if_link/if_choice_transition
      -- CP-element group 50: 	 branch_block_stmt_9401/if_stmt_9471_if_link/$exit
      -- 
    if_choice_transition_1281_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_9471_branch_ack_1, ack => Out_wrap_daemon_CP_855_elements(50)); -- 
    -- CP-element group 51:  transition  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	48 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	52 
    -- CP-element group 51:  members (1) 
      -- CP-element group 51: 	 branch_block_stmt_9401/if_stmt_9471_else_link/$entry
      -- 
    Out_wrap_daemon_CP_855_elements(51) <= Out_wrap_daemon_CP_855_elements(48);
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	51 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	54 
    -- CP-element group 52:  members (2) 
      -- CP-element group 52: 	 branch_block_stmt_9401/if_stmt_9471_else_link/$exit
      -- CP-element group 52: 	 branch_block_stmt_9401/if_stmt_9471_else_link/else_choice_transition
      -- 
    else_choice_transition_1285_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_9471_branch_ack_0, ack => Out_wrap_daemon_CP_855_elements(52)); -- 
    -- CP-element group 53:  place  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	50 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	96 
    -- CP-element group 53:  members (1) 
      -- CP-element group 53: 	 branch_block_stmt_9401/loop1
      -- 
    Out_wrap_daemon_CP_855_elements(53) <= Out_wrap_daemon_CP_855_elements(50);
    -- CP-element group 54:  branch  place  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	52 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	56 
    -- CP-element group 54: 	57 
    -- CP-element group 54:  members (1) 
      -- CP-element group 54: 	 branch_block_stmt_9401/if_stmt_9477__entry__
      -- 
    Out_wrap_daemon_CP_855_elements(54) <= Out_wrap_daemon_CP_855_elements(52);
    -- CP-element group 55:  merge  place  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	62 
    -- CP-element group 55: 	67 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	103 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 branch_block_stmt_9401/if_stmt_9477__exit__
      -- CP-element group 55: 	 branch_block_stmt_9401/branch_block_stmt_9401__exit__
      -- CP-element group 55: 	 branch_block_stmt_9401/if_stmt_9471__exit__
      -- 
    Out_wrap_daemon_CP_855_elements(55) <= OrReduce(Out_wrap_daemon_CP_855_elements(62) & Out_wrap_daemon_CP_855_elements(67));
    -- CP-element group 56:  transition  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	54 
    -- CP-element group 56: successors 
    -- CP-element group 56:  members (1) 
      -- CP-element group 56: 	 branch_block_stmt_9401/if_stmt_9477_dead_link/$entry
      -- 
    Out_wrap_daemon_CP_855_elements(56) <= Out_wrap_daemon_CP_855_elements(54);
    -- CP-element group 57:  transition  output  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	54 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57:  members (17) 
      -- CP-element group 57: 	 branch_block_stmt_9401/if_stmt_9477_eval_test/ULT_u15_u1_9480/ULT_u15_u1_9480_inputs/$entry
      -- CP-element group 57: 	 branch_block_stmt_9401/if_stmt_9477_eval_test/ULT_u15_u1_9480/ULT_u15_u1_9480_inputs/$exit
      -- CP-element group 57: 	 branch_block_stmt_9401/if_stmt_9477_eval_test/ULT_u15_u1_9480/SplitProtocol/Sample/rr
      -- CP-element group 57: 	 branch_block_stmt_9401/if_stmt_9477_eval_test/ULT_u15_u1_9480/SplitProtocol/Sample/$entry
      -- CP-element group 57: 	 branch_block_stmt_9401/if_stmt_9477_eval_test/ULT_u15_u1_9480/SplitProtocol/Sample/$exit
      -- CP-element group 57: 	 branch_block_stmt_9401/if_stmt_9477_eval_test/ULT_u15_u1_9480/SplitProtocol/$entry
      -- CP-element group 57: 	 branch_block_stmt_9401/if_stmt_9477_eval_test/ULT_u15_u1_9480/SplitProtocol/$exit
      -- CP-element group 57: 	 branch_block_stmt_9401/if_stmt_9477_eval_test/ULT_u15_u1_9480/$entry
      -- CP-element group 57: 	 branch_block_stmt_9401/if_stmt_9477_eval_test/ULT_u15_u1_9480/$exit
      -- CP-element group 57: 	 branch_block_stmt_9401/if_stmt_9477_eval_test/branch_req
      -- CP-element group 57: 	 branch_block_stmt_9401/if_stmt_9477_eval_test/$entry
      -- CP-element group 57: 	 branch_block_stmt_9401/if_stmt_9477_eval_test/ULT_u15_u1_9480/SplitProtocol/Update/cr
      -- CP-element group 57: 	 branch_block_stmt_9401/if_stmt_9477_eval_test/ULT_u15_u1_9480/SplitProtocol/Update/ca
      -- CP-element group 57: 	 branch_block_stmt_9401/if_stmt_9477_eval_test/ULT_u15_u1_9480/SplitProtocol/Update/$entry
      -- CP-element group 57: 	 branch_block_stmt_9401/if_stmt_9477_eval_test/ULT_u15_u1_9480/SplitProtocol/Update/$exit
      -- CP-element group 57: 	 branch_block_stmt_9401/if_stmt_9477_eval_test/$exit
      -- CP-element group 57: 	 branch_block_stmt_9401/if_stmt_9477_eval_test/ULT_u15_u1_9480/SplitProtocol/Sample/ra
      -- 
    branch_req_1315_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1315_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => Out_wrap_daemon_CP_855_elements(57), ack => if_stmt_9477_branch_req_0); -- 
    Out_wrap_daemon_CP_855_elements(57) <= Out_wrap_daemon_CP_855_elements(54);
    -- CP-element group 58:  branch  place  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	57 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58: 	61 
    -- CP-element group 58:  members (1) 
      -- CP-element group 58: 	 branch_block_stmt_9401/ULT_u15_u1_9480_place
      -- 
    Out_wrap_daemon_CP_855_elements(58) <= Out_wrap_daemon_CP_855_elements(57);
    -- CP-element group 59:  transition  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	60 
    -- CP-element group 59:  members (1) 
      -- CP-element group 59: 	 branch_block_stmt_9401/if_stmt_9477_if_link/$entry
      -- 
    Out_wrap_daemon_CP_855_elements(59) <= Out_wrap_daemon_CP_855_elements(58);
    -- CP-element group 60:  transition  input  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	59 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	63 
    -- CP-element group 60:  members (2) 
      -- CP-element group 60: 	 branch_block_stmt_9401/if_stmt_9477_if_link/$exit
      -- CP-element group 60: 	 branch_block_stmt_9401/if_stmt_9477_if_link/if_choice_transition
      -- 
    if_choice_transition_1320_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_9477_branch_ack_1, ack => Out_wrap_daemon_CP_855_elements(60)); -- 
    -- CP-element group 61:  transition  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	58 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	62 
    -- CP-element group 61:  members (1) 
      -- CP-element group 61: 	 branch_block_stmt_9401/if_stmt_9477_else_link/$entry
      -- 
    Out_wrap_daemon_CP_855_elements(61) <= Out_wrap_daemon_CP_855_elements(58);
    -- CP-element group 62:  transition  input  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	61 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	55 
    -- CP-element group 62:  members (2) 
      -- CP-element group 62: 	 branch_block_stmt_9401/if_stmt_9477_else_link/$exit
      -- CP-element group 62: 	 branch_block_stmt_9401/if_stmt_9477_else_link/else_choice_transition
      -- 
    else_choice_transition_1324_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_9477_branch_ack_0, ack => Out_wrap_daemon_CP_855_elements(62)); -- 
    -- CP-element group 63:  branch  place  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	60 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	82 
    -- CP-element group 63: 	83 
    -- CP-element group 63:  members (1) 
      -- CP-element group 63: 	 branch_block_stmt_9401/merge_stmt_9481__entry__
      -- 
    Out_wrap_daemon_CP_855_elements(63) <= Out_wrap_daemon_CP_855_elements(60);
    -- CP-element group 64:  merge  place  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	93 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	68 
    -- CP-element group 64:  members (2) 
      -- CP-element group 64: 	 branch_block_stmt_9401/assign_stmt_9489__entry__
      -- CP-element group 64: 	 branch_block_stmt_9401/merge_stmt_9481__exit__
      -- 
    Out_wrap_daemon_CP_855_elements(64) <= Out_wrap_daemon_CP_855_elements(93);
    -- CP-element group 65:  place  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	72 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	73 
    -- CP-element group 65:  members (2) 
      -- CP-element group 65: 	 branch_block_stmt_9401/assign_stmt_9494__entry__
      -- CP-element group 65: 	 branch_block_stmt_9401/assign_stmt_9489__exit__
      -- 
    Out_wrap_daemon_CP_855_elements(65) <= Out_wrap_daemon_CP_855_elements(72);
    -- CP-element group 66:  branch  place  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	73 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	74 
    -- CP-element group 66: 	75 
    -- CP-element group 66:  members (2) 
      -- CP-element group 66: 	 branch_block_stmt_9401/assign_stmt_9494__exit__
      -- CP-element group 66: 	 branch_block_stmt_9401/if_stmt_9495__entry__
      -- 
    Out_wrap_daemon_CP_855_elements(66) <= Out_wrap_daemon_CP_855_elements(73);
    -- CP-element group 67:  merge  place  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	80 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	55 
    -- CP-element group 67:  members (1) 
      -- CP-element group 67: 	 branch_block_stmt_9401/if_stmt_9495__exit__
      -- 
    Out_wrap_daemon_CP_855_elements(67) <= Out_wrap_daemon_CP_855_elements(80);
    -- CP-element group 68:  transition  output  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	64 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	69 
    -- CP-element group 68:  members (4) 
      -- CP-element group 68: 	 branch_block_stmt_9401/assign_stmt_9489/RPIPE_out_wrap_data_9488_Sample/rr
      -- CP-element group 68: 	 branch_block_stmt_9401/assign_stmt_9489/$entry
      -- CP-element group 68: 	 branch_block_stmt_9401/assign_stmt_9489/RPIPE_out_wrap_data_9488_sample_start_
      -- CP-element group 68: 	 branch_block_stmt_9401/assign_stmt_9489/RPIPE_out_wrap_data_9488_Sample/$entry
      -- 
    rr_1343_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1343_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => Out_wrap_daemon_CP_855_elements(68), ack => RPIPE_out_wrap_data_9488_inst_req_0); -- 
    Out_wrap_daemon_CP_855_elements(68) <= Out_wrap_daemon_CP_855_elements(64);
    -- CP-element group 69:  transition  input  output  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	68 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	70 
    -- CP-element group 69:  members (6) 
      -- CP-element group 69: 	 branch_block_stmt_9401/assign_stmt_9489/RPIPE_out_wrap_data_9488_Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_9401/assign_stmt_9489/RPIPE_out_wrap_data_9488_Update/cr
      -- CP-element group 69: 	 branch_block_stmt_9401/assign_stmt_9489/RPIPE_out_wrap_data_9488_Sample/ra
      -- CP-element group 69: 	 branch_block_stmt_9401/assign_stmt_9489/RPIPE_out_wrap_data_9488_Sample/$exit
      -- CP-element group 69: 	 branch_block_stmt_9401/assign_stmt_9489/RPIPE_out_wrap_data_9488_update_start_
      -- CP-element group 69: 	 branch_block_stmt_9401/assign_stmt_9489/RPIPE_out_wrap_data_9488_sample_completed_
      -- 
    ra_1344_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_out_wrap_data_9488_inst_ack_0, ack => Out_wrap_daemon_CP_855_elements(69)); -- 
    cr_1348_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1348_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => Out_wrap_daemon_CP_855_elements(69), ack => RPIPE_out_wrap_data_9488_inst_req_1); -- 
    -- CP-element group 70:  transition  input  output  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	69 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70:  members (6) 
      -- CP-element group 70: 	 branch_block_stmt_9401/assign_stmt_9489/RPIPE_out_wrap_data_9488_Update/ca
      -- CP-element group 70: 	 branch_block_stmt_9401/assign_stmt_9489/WPIPE_w_out_buf_9487_sample_start_
      -- CP-element group 70: 	 branch_block_stmt_9401/assign_stmt_9489/RPIPE_out_wrap_data_9488_update_completed_
      -- CP-element group 70: 	 branch_block_stmt_9401/assign_stmt_9489/RPIPE_out_wrap_data_9488_Update/$exit
      -- CP-element group 70: 	 branch_block_stmt_9401/assign_stmt_9489/WPIPE_w_out_buf_9487_Sample/req
      -- CP-element group 70: 	 branch_block_stmt_9401/assign_stmt_9489/WPIPE_w_out_buf_9487_Sample/$entry
      -- 
    ca_1349_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_out_wrap_data_9488_inst_ack_1, ack => Out_wrap_daemon_CP_855_elements(70)); -- 
    req_1357_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1357_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => Out_wrap_daemon_CP_855_elements(70), ack => WPIPE_w_out_buf_9487_inst_req_0); -- 
    -- CP-element group 71:  transition  input  output  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	72 
    -- CP-element group 71:  members (6) 
      -- CP-element group 71: 	 branch_block_stmt_9401/assign_stmt_9489/WPIPE_w_out_buf_9487_sample_completed_
      -- CP-element group 71: 	 branch_block_stmt_9401/assign_stmt_9489/WPIPE_w_out_buf_9487_update_start_
      -- CP-element group 71: 	 branch_block_stmt_9401/assign_stmt_9489/WPIPE_w_out_buf_9487_Sample/ack
      -- CP-element group 71: 	 branch_block_stmt_9401/assign_stmt_9489/WPIPE_w_out_buf_9487_Sample/$exit
      -- CP-element group 71: 	 branch_block_stmt_9401/assign_stmt_9489/WPIPE_w_out_buf_9487_Update/$entry
      -- CP-element group 71: 	 branch_block_stmt_9401/assign_stmt_9489/WPIPE_w_out_buf_9487_Update/req
      -- 
    ack_1358_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_w_out_buf_9487_inst_ack_0, ack => Out_wrap_daemon_CP_855_elements(71)); -- 
    req_1362_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1362_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => Out_wrap_daemon_CP_855_elements(71), ack => WPIPE_w_out_buf_9487_inst_req_1); -- 
    -- CP-element group 72:  transition  input  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	71 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	65 
    -- CP-element group 72:  members (4) 
      -- CP-element group 72: 	 branch_block_stmt_9401/assign_stmt_9489/$exit
      -- CP-element group 72: 	 branch_block_stmt_9401/assign_stmt_9489/WPIPE_w_out_buf_9487_update_completed_
      -- CP-element group 72: 	 branch_block_stmt_9401/assign_stmt_9489/WPIPE_w_out_buf_9487_Update/$exit
      -- CP-element group 72: 	 branch_block_stmt_9401/assign_stmt_9489/WPIPE_w_out_buf_9487_Update/ack
      -- 
    ack_1363_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_w_out_buf_9487_inst_ack_1, ack => Out_wrap_daemon_CP_855_elements(72)); -- 
    -- CP-element group 73:  transition  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	65 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	66 
    -- CP-element group 73:  members (18) 
      -- CP-element group 73: 	 branch_block_stmt_9401/assign_stmt_9494/$entry
      -- CP-element group 73: 	 branch_block_stmt_9401/assign_stmt_9494/$exit
      -- CP-element group 73: 	 branch_block_stmt_9401/assign_stmt_9494/ADD_u15_u15_9493_sample_start_
      -- CP-element group 73: 	 branch_block_stmt_9401/assign_stmt_9494/ADD_u15_u15_9493_sample_completed_
      -- CP-element group 73: 	 branch_block_stmt_9401/assign_stmt_9494/ADD_u15_u15_9493_update_start_
      -- CP-element group 73: 	 branch_block_stmt_9401/assign_stmt_9494/ADD_u15_u15_9493_update_completed_
      -- CP-element group 73: 	 branch_block_stmt_9401/assign_stmt_9494/R_count_var2_9491_sample_start_
      -- CP-element group 73: 	 branch_block_stmt_9401/assign_stmt_9494/R_count_var2_9491_sample_completed_
      -- CP-element group 73: 	 branch_block_stmt_9401/assign_stmt_9494/R_count_var2_9491_update_start_
      -- CP-element group 73: 	 branch_block_stmt_9401/assign_stmt_9494/R_count_var2_9491_update_completed_
      -- CP-element group 73: 	 branch_block_stmt_9401/assign_stmt_9494/ADD_u15_u15_9493_Sample/$entry
      -- CP-element group 73: 	 branch_block_stmt_9401/assign_stmt_9494/ADD_u15_u15_9493_Sample/$exit
      -- CP-element group 73: 	 branch_block_stmt_9401/assign_stmt_9494/ADD_u15_u15_9493_Sample/rr
      -- CP-element group 73: 	 branch_block_stmt_9401/assign_stmt_9494/ADD_u15_u15_9493_Sample/ra
      -- CP-element group 73: 	 branch_block_stmt_9401/assign_stmt_9494/ADD_u15_u15_9493_Update/$entry
      -- CP-element group 73: 	 branch_block_stmt_9401/assign_stmt_9494/ADD_u15_u15_9493_Update/$exit
      -- CP-element group 73: 	 branch_block_stmt_9401/assign_stmt_9494/ADD_u15_u15_9493_Update/cr
      -- CP-element group 73: 	 branch_block_stmt_9401/assign_stmt_9494/ADD_u15_u15_9493_Update/ca
      -- 
    Out_wrap_daemon_CP_855_elements(73) <= Out_wrap_daemon_CP_855_elements(65);
    -- CP-element group 74:  transition  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	66 
    -- CP-element group 74: successors 
    -- CP-element group 74:  members (1) 
      -- CP-element group 74: 	 branch_block_stmt_9401/if_stmt_9495_dead_link/$entry
      -- 
    Out_wrap_daemon_CP_855_elements(74) <= Out_wrap_daemon_CP_855_elements(66);
    -- CP-element group 75:  transition  output  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	66 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	76 
    -- CP-element group 75:  members (17) 
      -- CP-element group 75: 	 branch_block_stmt_9401/if_stmt_9495_eval_test/$entry
      -- CP-element group 75: 	 branch_block_stmt_9401/if_stmt_9495_eval_test/$exit
      -- CP-element group 75: 	 branch_block_stmt_9401/if_stmt_9495_eval_test/ULT_u15_u1_9498/$entry
      -- CP-element group 75: 	 branch_block_stmt_9401/if_stmt_9495_eval_test/ULT_u15_u1_9498/$exit
      -- CP-element group 75: 	 branch_block_stmt_9401/if_stmt_9495_eval_test/ULT_u15_u1_9498/ULT_u15_u1_9498_inputs/$entry
      -- CP-element group 75: 	 branch_block_stmt_9401/if_stmt_9495_eval_test/ULT_u15_u1_9498/ULT_u15_u1_9498_inputs/$exit
      -- CP-element group 75: 	 branch_block_stmt_9401/if_stmt_9495_eval_test/ULT_u15_u1_9498/SplitProtocol/$entry
      -- CP-element group 75: 	 branch_block_stmt_9401/if_stmt_9495_eval_test/ULT_u15_u1_9498/SplitProtocol/$exit
      -- CP-element group 75: 	 branch_block_stmt_9401/if_stmt_9495_eval_test/ULT_u15_u1_9498/SplitProtocol/Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_9401/if_stmt_9495_eval_test/ULT_u15_u1_9498/SplitProtocol/Sample/$exit
      -- CP-element group 75: 	 branch_block_stmt_9401/if_stmt_9495_eval_test/ULT_u15_u1_9498/SplitProtocol/Sample/rr
      -- CP-element group 75: 	 branch_block_stmt_9401/if_stmt_9495_eval_test/ULT_u15_u1_9498/SplitProtocol/Sample/ra
      -- CP-element group 75: 	 branch_block_stmt_9401/if_stmt_9495_eval_test/ULT_u15_u1_9498/SplitProtocol/Update/$entry
      -- CP-element group 75: 	 branch_block_stmt_9401/if_stmt_9495_eval_test/ULT_u15_u1_9498/SplitProtocol/Update/$exit
      -- CP-element group 75: 	 branch_block_stmt_9401/if_stmt_9495_eval_test/ULT_u15_u1_9498/SplitProtocol/Update/cr
      -- CP-element group 75: 	 branch_block_stmt_9401/if_stmt_9495_eval_test/ULT_u15_u1_9498/SplitProtocol/Update/ca
      -- CP-element group 75: 	 branch_block_stmt_9401/if_stmt_9495_eval_test/branch_req
      -- 
    branch_req_1411_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1411_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => Out_wrap_daemon_CP_855_elements(75), ack => if_stmt_9495_branch_req_0); -- 
    Out_wrap_daemon_CP_855_elements(75) <= Out_wrap_daemon_CP_855_elements(66);
    -- CP-element group 76:  branch  place  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	75 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	77 
    -- CP-element group 76: 	79 
    -- CP-element group 76:  members (1) 
      -- CP-element group 76: 	 branch_block_stmt_9401/ULT_u15_u1_9498_place
      -- 
    Out_wrap_daemon_CP_855_elements(76) <= Out_wrap_daemon_CP_855_elements(75);
    -- CP-element group 77:  transition  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	76 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	78 
    -- CP-element group 77:  members (1) 
      -- CP-element group 77: 	 branch_block_stmt_9401/if_stmt_9495_if_link/$entry
      -- 
    Out_wrap_daemon_CP_855_elements(77) <= Out_wrap_daemon_CP_855_elements(76);
    -- CP-element group 78:  transition  input  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	77 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	81 
    -- CP-element group 78:  members (2) 
      -- CP-element group 78: 	 branch_block_stmt_9401/if_stmt_9495_if_link/$exit
      -- CP-element group 78: 	 branch_block_stmt_9401/if_stmt_9495_if_link/if_choice_transition
      -- 
    if_choice_transition_1416_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_9495_branch_ack_1, ack => Out_wrap_daemon_CP_855_elements(78)); -- 
    -- CP-element group 79:  transition  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	76 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	80 
    -- CP-element group 79:  members (1) 
      -- CP-element group 79: 	 branch_block_stmt_9401/if_stmt_9495_else_link/$entry
      -- 
    Out_wrap_daemon_CP_855_elements(79) <= Out_wrap_daemon_CP_855_elements(76);
    -- CP-element group 80:  transition  input  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	79 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	67 
    -- CP-element group 80:  members (2) 
      -- CP-element group 80: 	 branch_block_stmt_9401/if_stmt_9495_else_link/$exit
      -- CP-element group 80: 	 branch_block_stmt_9401/if_stmt_9495_else_link/else_choice_transition
      -- 
    else_choice_transition_1420_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_9495_branch_ack_0, ack => Out_wrap_daemon_CP_855_elements(80)); -- 
    -- CP-element group 81:  place  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	78 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	87 
    -- CP-element group 81:  members (1) 
      -- CP-element group 81: 	 branch_block_stmt_9401/loop2
      -- 
    Out_wrap_daemon_CP_855_elements(81) <= Out_wrap_daemon_CP_855_elements(78);
    -- CP-element group 82:  transition  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	63 
    -- CP-element group 82: successors 
    -- CP-element group 82:  members (1) 
      -- CP-element group 82: 	 branch_block_stmt_9401/merge_stmt_9481_dead_link/$entry
      -- 
    Out_wrap_daemon_CP_855_elements(82) <= Out_wrap_daemon_CP_855_elements(63);
    -- CP-element group 83:  fork  transition  output  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	63 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	84 
    -- CP-element group 83: 	85 
    -- CP-element group 83:  members (8) 
      -- CP-element group 83: 	 branch_block_stmt_9401/merge_stmt_9481__entry___PhiReq/$entry
      -- CP-element group 83: 	 branch_block_stmt_9401/merge_stmt_9481__entry___PhiReq/phi_stmt_9482/$entry
      -- CP-element group 83: 	 branch_block_stmt_9401/merge_stmt_9481__entry___PhiReq/phi_stmt_9482/phi_stmt_9482_sources/$entry
      -- CP-element group 83: 	 branch_block_stmt_9401/merge_stmt_9481__entry___PhiReq/phi_stmt_9482/phi_stmt_9482_sources/Interlock/$entry
      -- CP-element group 83: 	 branch_block_stmt_9401/merge_stmt_9481__entry___PhiReq/phi_stmt_9482/phi_stmt_9482_sources/Interlock/Sample/$entry
      -- CP-element group 83: 	 branch_block_stmt_9401/merge_stmt_9481__entry___PhiReq/phi_stmt_9482/phi_stmt_9482_sources/Interlock/Sample/req
      -- CP-element group 83: 	 branch_block_stmt_9401/merge_stmt_9481__entry___PhiReq/phi_stmt_9482/phi_stmt_9482_sources/Interlock/Update/$entry
      -- CP-element group 83: 	 branch_block_stmt_9401/merge_stmt_9481__entry___PhiReq/phi_stmt_9482/phi_stmt_9482_sources/Interlock/Update/req
      -- 
    req_1441_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1441_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => Out_wrap_daemon_CP_855_elements(83), ack => n_count_var_9470_9484_buf_req_0); -- 
    req_1446_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1446_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => Out_wrap_daemon_CP_855_elements(83), ack => n_count_var_9470_9484_buf_req_1); -- 
    Out_wrap_daemon_CP_855_elements(83) <= Out_wrap_daemon_CP_855_elements(63);
    -- CP-element group 84:  transition  input  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	83 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	86 
    -- CP-element group 84:  members (2) 
      -- CP-element group 84: 	 branch_block_stmt_9401/merge_stmt_9481__entry___PhiReq/phi_stmt_9482/phi_stmt_9482_sources/Interlock/Sample/$exit
      -- CP-element group 84: 	 branch_block_stmt_9401/merge_stmt_9481__entry___PhiReq/phi_stmt_9482/phi_stmt_9482_sources/Interlock/Sample/ack
      -- 
    ack_1442_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_count_var_9470_9484_buf_ack_0, ack => Out_wrap_daemon_CP_855_elements(84)); -- 
    -- CP-element group 85:  transition  input  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	83 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	86 
    -- CP-element group 85:  members (2) 
      -- CP-element group 85: 	 branch_block_stmt_9401/merge_stmt_9481__entry___PhiReq/phi_stmt_9482/phi_stmt_9482_sources/Interlock/Update/$exit
      -- CP-element group 85: 	 branch_block_stmt_9401/merge_stmt_9481__entry___PhiReq/phi_stmt_9482/phi_stmt_9482_sources/Interlock/Update/ack
      -- 
    ack_1447_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_count_var_9470_9484_buf_ack_1, ack => Out_wrap_daemon_CP_855_elements(85)); -- 
    -- CP-element group 86:  join  transition  output  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	84 
    -- CP-element group 86: 	85 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	91 
    -- CP-element group 86:  members (5) 
      -- CP-element group 86: 	 branch_block_stmt_9401/merge_stmt_9481__entry___PhiReq/$exit
      -- CP-element group 86: 	 branch_block_stmt_9401/merge_stmt_9481__entry___PhiReq/phi_stmt_9482/$exit
      -- CP-element group 86: 	 branch_block_stmt_9401/merge_stmt_9481__entry___PhiReq/phi_stmt_9482/phi_stmt_9482_sources/$exit
      -- CP-element group 86: 	 branch_block_stmt_9401/merge_stmt_9481__entry___PhiReq/phi_stmt_9482/phi_stmt_9482_sources/Interlock/$exit
      -- CP-element group 86: 	 branch_block_stmt_9401/merge_stmt_9481__entry___PhiReq/phi_stmt_9482/phi_stmt_9482_req
      -- 
    phi_stmt_9482_req_1448_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_9482_req_1448_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => Out_wrap_daemon_CP_855_elements(86), ack => phi_stmt_9482_req_0); -- 
    Out_wrap_daemon_cp_element_group_86: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "Out_wrap_daemon_cp_element_group_86"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= Out_wrap_daemon_CP_855_elements(84) & Out_wrap_daemon_CP_855_elements(85);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => Out_wrap_daemon_CP_855_elements(86), clk => clk, reset => reset); --
    end block;
    -- CP-element group 87:  fork  transition  output  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	81 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87: 	89 
    -- CP-element group 87:  members (8) 
      -- CP-element group 87: 	 branch_block_stmt_9401/loop2_PhiReq/$entry
      -- CP-element group 87: 	 branch_block_stmt_9401/loop2_PhiReq/phi_stmt_9482/$entry
      -- CP-element group 87: 	 branch_block_stmt_9401/loop2_PhiReq/phi_stmt_9482/phi_stmt_9482_sources/$entry
      -- CP-element group 87: 	 branch_block_stmt_9401/loop2_PhiReq/phi_stmt_9482/phi_stmt_9482_sources/Interlock/$entry
      -- CP-element group 87: 	 branch_block_stmt_9401/loop2_PhiReq/phi_stmt_9482/phi_stmt_9482_sources/Interlock/Sample/$entry
      -- CP-element group 87: 	 branch_block_stmt_9401/loop2_PhiReq/phi_stmt_9482/phi_stmt_9482_sources/Interlock/Sample/req
      -- CP-element group 87: 	 branch_block_stmt_9401/loop2_PhiReq/phi_stmt_9482/phi_stmt_9482_sources/Interlock/Update/$entry
      -- CP-element group 87: 	 branch_block_stmt_9401/loop2_PhiReq/phi_stmt_9482/phi_stmt_9482_sources/Interlock/Update/req
      -- 
    req_1464_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1464_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => Out_wrap_daemon_CP_855_elements(87), ack => n_count_var2_9494_9485_buf_req_0); -- 
    req_1469_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1469_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => Out_wrap_daemon_CP_855_elements(87), ack => n_count_var2_9494_9485_buf_req_1); -- 
    Out_wrap_daemon_CP_855_elements(87) <= Out_wrap_daemon_CP_855_elements(81);
    -- CP-element group 88:  transition  input  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	87 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	90 
    -- CP-element group 88:  members (2) 
      -- CP-element group 88: 	 branch_block_stmt_9401/loop2_PhiReq/phi_stmt_9482/phi_stmt_9482_sources/Interlock/Sample/$exit
      -- CP-element group 88: 	 branch_block_stmt_9401/loop2_PhiReq/phi_stmt_9482/phi_stmt_9482_sources/Interlock/Sample/ack
      -- 
    ack_1465_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_count_var2_9494_9485_buf_ack_0, ack => Out_wrap_daemon_CP_855_elements(88)); -- 
    -- CP-element group 89:  transition  input  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	87 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	90 
    -- CP-element group 89:  members (2) 
      -- CP-element group 89: 	 branch_block_stmt_9401/loop2_PhiReq/phi_stmt_9482/phi_stmt_9482_sources/Interlock/Update/$exit
      -- CP-element group 89: 	 branch_block_stmt_9401/loop2_PhiReq/phi_stmt_9482/phi_stmt_9482_sources/Interlock/Update/ack
      -- 
    ack_1470_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_count_var2_9494_9485_buf_ack_1, ack => Out_wrap_daemon_CP_855_elements(89)); -- 
    -- CP-element group 90:  join  transition  output  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	88 
    -- CP-element group 90: 	89 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	91 
    -- CP-element group 90:  members (5) 
      -- CP-element group 90: 	 branch_block_stmt_9401/loop2_PhiReq/$exit
      -- CP-element group 90: 	 branch_block_stmt_9401/loop2_PhiReq/phi_stmt_9482/$exit
      -- CP-element group 90: 	 branch_block_stmt_9401/loop2_PhiReq/phi_stmt_9482/phi_stmt_9482_sources/$exit
      -- CP-element group 90: 	 branch_block_stmt_9401/loop2_PhiReq/phi_stmt_9482/phi_stmt_9482_sources/Interlock/$exit
      -- CP-element group 90: 	 branch_block_stmt_9401/loop2_PhiReq/phi_stmt_9482/phi_stmt_9482_req
      -- 
    phi_stmt_9482_req_1471_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_9482_req_1471_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => Out_wrap_daemon_CP_855_elements(90), ack => phi_stmt_9482_req_1); -- 
    Out_wrap_daemon_cp_element_group_90: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "Out_wrap_daemon_cp_element_group_90"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= Out_wrap_daemon_CP_855_elements(88) & Out_wrap_daemon_CP_855_elements(89);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => Out_wrap_daemon_CP_855_elements(90), clk => clk, reset => reset); --
    end block;
    -- CP-element group 91:  merge  place  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	86 
    -- CP-element group 91: 	90 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	92 
    -- CP-element group 91:  members (1) 
      -- CP-element group 91: 	 branch_block_stmt_9401/merge_stmt_9481_PhiReqMerge
      -- 
    Out_wrap_daemon_CP_855_elements(91) <= OrReduce(Out_wrap_daemon_CP_855_elements(86) & Out_wrap_daemon_CP_855_elements(90));
    -- CP-element group 92:  transition  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	91 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	93 
    -- CP-element group 92:  members (1) 
      -- CP-element group 92: 	 branch_block_stmt_9401/merge_stmt_9481_PhiAck/$entry
      -- 
    Out_wrap_daemon_CP_855_elements(92) <= Out_wrap_daemon_CP_855_elements(91);
    -- CP-element group 93:  transition  input  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	92 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	64 
    -- CP-element group 93:  members (2) 
      -- CP-element group 93: 	 branch_block_stmt_9401/merge_stmt_9481_PhiAck/$exit
      -- CP-element group 93: 	 branch_block_stmt_9401/merge_stmt_9481_PhiAck/phi_stmt_9482_ack
      -- 
    phi_stmt_9482_ack_1476_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_9482_ack_0, ack => Out_wrap_daemon_CP_855_elements(93)); -- 
    -- CP-element group 94:  transition  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	5 
    -- CP-element group 94: successors 
    -- CP-element group 94:  members (1) 
      -- CP-element group 94: 	 branch_block_stmt_9401/merge_stmt_9448_dead_link/$entry
      -- 
    Out_wrap_daemon_CP_855_elements(94) <= Out_wrap_daemon_CP_855_elements(5);
    -- CP-element group 95:  transition  output  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	5 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	100 
    -- CP-element group 95:  members (7) 
      -- CP-element group 95: 	 branch_block_stmt_9401/merge_stmt_9448__entry___PhiReq/$entry
      -- CP-element group 95: 	 branch_block_stmt_9401/merge_stmt_9448__entry___PhiReq/$exit
      -- CP-element group 95: 	 branch_block_stmt_9401/merge_stmt_9448__entry___PhiReq/phi_stmt_9449/$entry
      -- CP-element group 95: 	 branch_block_stmt_9401/merge_stmt_9448__entry___PhiReq/phi_stmt_9449/$exit
      -- CP-element group 95: 	 branch_block_stmt_9401/merge_stmt_9448__entry___PhiReq/phi_stmt_9449/phi_stmt_9449_sources/$entry
      -- CP-element group 95: 	 branch_block_stmt_9401/merge_stmt_9448__entry___PhiReq/phi_stmt_9449/phi_stmt_9449_sources/$exit
      -- CP-element group 95: 	 branch_block_stmt_9401/merge_stmt_9448__entry___PhiReq/phi_stmt_9449/phi_stmt_9449_req
      -- 
    phi_stmt_9449_req_1490_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_9449_req_1490_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => Out_wrap_daemon_CP_855_elements(95), ack => phi_stmt_9449_req_0); -- 
    Out_wrap_daemon_CP_855_elements(95) <= Out_wrap_daemon_CP_855_elements(5);
    -- CP-element group 96:  fork  transition  output  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	53 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	97 
    -- CP-element group 96: 	98 
    -- CP-element group 96:  members (8) 
      -- CP-element group 96: 	 branch_block_stmt_9401/loop1_PhiReq/$entry
      -- CP-element group 96: 	 branch_block_stmt_9401/loop1_PhiReq/phi_stmt_9449/$entry
      -- CP-element group 96: 	 branch_block_stmt_9401/loop1_PhiReq/phi_stmt_9449/phi_stmt_9449_sources/$entry
      -- CP-element group 96: 	 branch_block_stmt_9401/loop1_PhiReq/phi_stmt_9449/phi_stmt_9449_sources/Interlock/$entry
      -- CP-element group 96: 	 branch_block_stmt_9401/loop1_PhiReq/phi_stmt_9449/phi_stmt_9449_sources/Interlock/Sample/$entry
      -- CP-element group 96: 	 branch_block_stmt_9401/loop1_PhiReq/phi_stmt_9449/phi_stmt_9449_sources/Interlock/Sample/req
      -- CP-element group 96: 	 branch_block_stmt_9401/loop1_PhiReq/phi_stmt_9449/phi_stmt_9449_sources/Interlock/Update/$entry
      -- CP-element group 96: 	 branch_block_stmt_9401/loop1_PhiReq/phi_stmt_9449/phi_stmt_9449_sources/Interlock/Update/req
      -- 
    req_1506_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1506_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => Out_wrap_daemon_CP_855_elements(96), ack => n_count_var_9470_9452_buf_req_0); -- 
    req_1511_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1511_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => Out_wrap_daemon_CP_855_elements(96), ack => n_count_var_9470_9452_buf_req_1); -- 
    Out_wrap_daemon_CP_855_elements(96) <= Out_wrap_daemon_CP_855_elements(53);
    -- CP-element group 97:  transition  input  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	96 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	99 
    -- CP-element group 97:  members (2) 
      -- CP-element group 97: 	 branch_block_stmt_9401/loop1_PhiReq/phi_stmt_9449/phi_stmt_9449_sources/Interlock/Sample/$exit
      -- CP-element group 97: 	 branch_block_stmt_9401/loop1_PhiReq/phi_stmt_9449/phi_stmt_9449_sources/Interlock/Sample/ack
      -- 
    ack_1507_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_count_var_9470_9452_buf_ack_0, ack => Out_wrap_daemon_CP_855_elements(97)); -- 
    -- CP-element group 98:  transition  input  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	96 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	99 
    -- CP-element group 98:  members (2) 
      -- CP-element group 98: 	 branch_block_stmt_9401/loop1_PhiReq/phi_stmt_9449/phi_stmt_9449_sources/Interlock/Update/$exit
      -- CP-element group 98: 	 branch_block_stmt_9401/loop1_PhiReq/phi_stmt_9449/phi_stmt_9449_sources/Interlock/Update/ack
      -- 
    ack_1512_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_count_var_9470_9452_buf_ack_1, ack => Out_wrap_daemon_CP_855_elements(98)); -- 
    -- CP-element group 99:  join  transition  output  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	97 
    -- CP-element group 99: 	98 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	100 
    -- CP-element group 99:  members (5) 
      -- CP-element group 99: 	 branch_block_stmt_9401/loop1_PhiReq/$exit
      -- CP-element group 99: 	 branch_block_stmt_9401/loop1_PhiReq/phi_stmt_9449/$exit
      -- CP-element group 99: 	 branch_block_stmt_9401/loop1_PhiReq/phi_stmt_9449/phi_stmt_9449_sources/$exit
      -- CP-element group 99: 	 branch_block_stmt_9401/loop1_PhiReq/phi_stmt_9449/phi_stmt_9449_sources/Interlock/$exit
      -- CP-element group 99: 	 branch_block_stmt_9401/loop1_PhiReq/phi_stmt_9449/phi_stmt_9449_req
      -- 
    phi_stmt_9449_req_1513_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_9449_req_1513_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => Out_wrap_daemon_CP_855_elements(99), ack => phi_stmt_9449_req_1); -- 
    Out_wrap_daemon_cp_element_group_99: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "Out_wrap_daemon_cp_element_group_99"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= Out_wrap_daemon_CP_855_elements(97) & Out_wrap_daemon_CP_855_elements(98);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => Out_wrap_daemon_CP_855_elements(99), clk => clk, reset => reset); --
    end block;
    -- CP-element group 100:  merge  place  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	95 
    -- CP-element group 100: 	99 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	101 
    -- CP-element group 100:  members (1) 
      -- CP-element group 100: 	 branch_block_stmt_9401/merge_stmt_9448_PhiReqMerge
      -- 
    Out_wrap_daemon_CP_855_elements(100) <= OrReduce(Out_wrap_daemon_CP_855_elements(95) & Out_wrap_daemon_CP_855_elements(99));
    -- CP-element group 101:  transition  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	100 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	102 
    -- CP-element group 101:  members (1) 
      -- CP-element group 101: 	 branch_block_stmt_9401/merge_stmt_9448_PhiAck/$entry
      -- 
    Out_wrap_daemon_CP_855_elements(101) <= Out_wrap_daemon_CP_855_elements(100);
    -- CP-element group 102:  transition  input  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	101 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	6 
    -- CP-element group 102:  members (2) 
      -- CP-element group 102: 	 branch_block_stmt_9401/merge_stmt_9448_PhiAck/$exit
      -- CP-element group 102: 	 branch_block_stmt_9401/merge_stmt_9448_PhiAck/phi_stmt_9449_ack
      -- 
    phi_stmt_9449_ack_1518_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_9449_ack_0, ack => Out_wrap_daemon_CP_855_elements(102)); -- 
    -- CP-element group 103:  transition  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	55 
    -- CP-element group 103: successors 
    -- CP-element group 103:  members (2) 
      -- CP-element group 103: 	 $exit
      -- CP-element group 103: 	 branch_block_stmt_9401/$exit
      -- 
    Out_wrap_daemon_CP_855_elements(103) <= Out_wrap_daemon_CP_855_elements(55);
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal CONCAT_u64_u128_9411_wire : std_logic_vector(127 downto 0);
    signal ED_9416 : std_logic_vector(0 downto 0);
    signal EQ_u1_u1_9457_wire : std_logic_vector(0 downto 0);
    signal MUX_9439_wire : std_logic_vector(14 downto 0);
    signal MUX_9445_wire : std_logic_vector(14 downto 0);
    signal RPIPE_d_out_buf_9463_wire : std_logic_vector(127 downto 0);
    signal RPIPE_e_out_buf_9459_wire : std_logic_vector(127 downto 0);
    signal RPIPE_out_wrap_data_9488_wire : std_logic_vector(127 downto 0);
    signal R_MAX_COUNT_9434_wire_constant : std_logic_vector(14 downto 0);
    signal R_MAX_COUNT_9437_wire_constant : std_logic_vector(14 downto 0);
    signal R_MAX_COUNT_9440_wire_constant : std_logic_vector(14 downto 0);
    signal R_MAX_COUNT_9479_wire_constant : std_logic_vector(14 downto 0);
    signal R_MAX_COUNT_9497_wire_constant : std_logic_vector(14 downto 0);
    signal R_ONE_COUNT_9451_wire_constant : std_logic_vector(14 downto 0);
    signal UGE_u15_u1_9442_wire : std_logic_vector(0 downto 0);
    signal ULT_u15_u1_9436_wire : std_logic_vector(0 downto 0);
    signal ULT_u15_u1_9474_wire : std_logic_vector(0 downto 0);
    signal ULT_u15_u1_9480_wire : std_logic_vector(0 downto 0);
    signal ULT_u15_u1_9498_wire : std_logic_vector(0 downto 0);
    signal count_9432 : std_logic_vector(14 downto 0);
    signal count_blocks_9447 : std_logic_vector(14 downto 0);
    signal count_var2_9482 : std_logic_vector(14 downto 0);
    signal count_var_9449 : std_logic_vector(14 downto 0);
    signal got_new_key_9424 : std_logic_vector(0 downto 0);
    signal head_out_9404 : std_logic_vector(63 downto 0);
    signal konst_9438_wire_constant : std_logic_vector(14 downto 0);
    signal konst_9444_wire_constant : std_logic_vector(14 downto 0);
    signal konst_9456_wire_constant : std_logic_vector(0 downto 0);
    signal konst_9468_wire_constant : std_logic_vector(14 downto 0);
    signal konst_9492_wire_constant : std_logic_vector(14 downto 0);
    signal mode_9420 : std_logic_vector(2 downto 0);
    signal n_count_var2_9494 : std_logic_vector(14 downto 0);
    signal n_count_var2_9494_9485_buffered : std_logic_vector(14 downto 0);
    signal n_count_var_9470 : std_logic_vector(14 downto 0);
    signal n_count_var_9470_9452_buffered : std_logic_vector(14 downto 0);
    signal n_count_var_9470_9484_buffered : std_logic_vector(14 downto 0);
    signal st_out_9407 : std_logic_vector(63 downto 0);
    signal unused_44_9428 : std_logic_vector(43 downto 0);
    signal xxOut_wrap_daemonxxMAX_COUNT : std_logic_vector(14 downto 0);
    signal xxOut_wrap_daemonxxONE_COUNT : std_logic_vector(14 downto 0);
    signal xxOut_wrap_daemonxxZERO : std_logic_vector(63 downto 0);
    signal xxOut_wrap_daemonxxZERO_COUNT : std_logic_vector(14 downto 0);
    -- 
  begin -- 
    R_MAX_COUNT_9434_wire_constant <= "000000111111111";
    R_MAX_COUNT_9437_wire_constant <= "000000111111111";
    R_MAX_COUNT_9440_wire_constant <= "000000111111111";
    R_MAX_COUNT_9479_wire_constant <= "000000111111111";
    R_MAX_COUNT_9497_wire_constant <= "000000111111111";
    R_ONE_COUNT_9451_wire_constant <= "000000000000001";
    konst_9438_wire_constant <= "000000000000000";
    konst_9444_wire_constant <= "000000000000000";
    konst_9456_wire_constant <= "0";
    konst_9468_wire_constant <= "000000000000001";
    konst_9492_wire_constant <= "000000000000001";
    xxOut_wrap_daemonxxMAX_COUNT <= "000000111111111";
    xxOut_wrap_daemonxxONE_COUNT <= "000000000000001";
    xxOut_wrap_daemonxxZERO <= "0000000000000000000000000000000000000000000000000000000000000000";
    xxOut_wrap_daemonxxZERO_COUNT <= "000000000000000";
    phi_stmt_9449: Block -- phi operator 
      signal idata: std_logic_vector(29 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ONE_COUNT_9451_wire_constant & n_count_var_9470_9452_buffered;
      req <= phi_stmt_9449_req_0 & phi_stmt_9449_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_9449",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 15) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_9449_ack_0,
          idata => idata,
          odata => count_var_9449,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_9449
    phi_stmt_9482: Block -- phi operator 
      signal idata: std_logic_vector(29 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= n_count_var_9470_9484_buffered & n_count_var2_9494_9485_buffered;
      req <= phi_stmt_9482_req_0 & phi_stmt_9482_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_9482",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 15) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_9482_ack_0,
          idata => idata,
          odata => count_var2_9482,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_9482
    -- flow-through select operator MUX_9439_inst
    MUX_9439_wire <= R_MAX_COUNT_9437_wire_constant when (ULT_u15_u1_9436_wire(0) /=  '0') else konst_9438_wire_constant;
    -- flow-through select operator MUX_9445_inst
    MUX_9445_wire <= count_9432 when (UGE_u15_u1_9442_wire(0) /=  '0') else konst_9444_wire_constant;
    -- flow-through slice operator slice_9415_inst
    ED_9416 <= head_out_9404(63 downto 63);
    -- flow-through slice operator slice_9419_inst
    mode_9420 <= head_out_9404(62 downto 60);
    -- flow-through slice operator slice_9423_inst
    got_new_key_9424 <= head_out_9404(59 downto 59);
    -- flow-through slice operator slice_9427_inst
    unused_44_9428 <= head_out_9404(58 downto 15);
    -- flow-through slice operator slice_9431_inst
    count_9432 <= head_out_9404(14 downto 0);
    n_count_var2_9494_9485_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_count_var2_9494_9485_buf_req_0;
      n_count_var2_9494_9485_buf_ack_0<= wack(0);
      rreq(0) <= n_count_var2_9494_9485_buf_req_1;
      n_count_var2_9494_9485_buf_ack_1<= rack(0);
      n_count_var2_9494_9485_buf : InterlockBuffer generic map ( -- 
        name => "n_count_var2_9494_9485_buf",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 15,
        out_data_width => 15,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_count_var2_9494,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_count_var2_9494_9485_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_count_var_9470_9452_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_count_var_9470_9452_buf_req_0;
      n_count_var_9470_9452_buf_ack_0<= wack(0);
      rreq(0) <= n_count_var_9470_9452_buf_req_1;
      n_count_var_9470_9452_buf_ack_1<= rack(0);
      n_count_var_9470_9452_buf : InterlockBuffer generic map ( -- 
        name => "n_count_var_9470_9452_buf",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 15,
        out_data_width => 15,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_count_var_9470,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_count_var_9470_9452_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_count_var_9470_9484_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_count_var_9470_9484_buf_req_0;
      n_count_var_9470_9484_buf_ack_0<= wack(0);
      rreq(0) <= n_count_var_9470_9484_buf_req_1;
      n_count_var_9470_9484_buf_ack_1<= rack(0);
      n_count_var_9470_9484_buf : InterlockBuffer generic map ( -- 
        name => "n_count_var_9470_9484_buf",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 15,
        out_data_width => 15,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_count_var_9470,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_count_var_9470_9484_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    if_stmt_9454_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= EQ_u1_u1_9457_wire;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_9454_branch", condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_9454_branch_req_0,
          ack0 => if_stmt_9454_branch_ack_0,
          ack1 => if_stmt_9454_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_9471_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= ULT_u15_u1_9474_wire;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_9471_branch", condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_9471_branch_req_0,
          ack0 => if_stmt_9471_branch_ack_0,
          ack1 => if_stmt_9471_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_9477_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= ULT_u15_u1_9480_wire;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_9477_branch", condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_9477_branch_req_0,
          ack0 => if_stmt_9477_branch_ack_0,
          ack1 => if_stmt_9477_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_9495_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= ULT_u15_u1_9498_wire;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_9495_branch", condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_9495_branch_req_0,
          ack0 => if_stmt_9495_branch_ack_0,
          ack1 => if_stmt_9495_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u15_u15_9469_inst
    process(count_var_9449) -- 
      variable tmp_var : std_logic_vector(14 downto 0); -- 
    begin -- 
      ApIntAdd_proc(count_var_9449, konst_9468_wire_constant, tmp_var);
      n_count_var_9470 <= tmp_var; -- 
    end process;
    -- binary operator ADD_u15_u15_9493_inst
    process(count_var2_9482) -- 
      variable tmp_var : std_logic_vector(14 downto 0); -- 
    begin -- 
      ApIntAdd_proc(count_var2_9482, konst_9492_wire_constant, tmp_var);
      n_count_var2_9494 <= tmp_var; -- 
    end process;
    -- shared split operator group (2) : CONCAT_u64_u128_9411_inst 
    ApConcat_group_2: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= head_out_9404 & st_out_9407;
      CONCAT_u64_u128_9411_wire <= data_out(127 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= CONCAT_u64_u128_9411_inst_req_0;
      CONCAT_u64_u128_9411_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= CONCAT_u64_u128_9411_inst_req_1;
      CONCAT_u64_u128_9411_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(name => "gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApConcat",
          name => "ApConcat_group_2",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 64, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 128,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 2
    -- binary operator EQ_u1_u1_9457_inst
    process(ED_9416) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(ED_9416, konst_9456_wire_constant, tmp_var);
      EQ_u1_u1_9457_wire <= tmp_var; -- 
    end process;
    -- shared split operator group (4) : OR_u15_u15_9446_inst 
    ApIntOr_group_4: Block -- 
      signal data_in: std_logic_vector(29 downto 0);
      signal data_out: std_logic_vector(14 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= MUX_9439_wire & MUX_9445_wire;
      count_blocks_9447 <= data_out(14 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= OR_u15_u15_9446_inst_req_0;
      OR_u15_u15_9446_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= OR_u15_u15_9446_inst_req_1;
      OR_u15_u15_9446_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(name => "gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          name => "ApIntOr_group_4",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 15,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 15, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 15,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 4
    -- binary operator UGE_u15_u1_9442_inst
    process(R_MAX_COUNT_9440_wire_constant, count_9432) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUge_proc(R_MAX_COUNT_9440_wire_constant, count_9432, tmp_var);
      UGE_u15_u1_9442_wire <= tmp_var; -- 
    end process;
    -- binary operator ULT_u15_u1_9436_inst
    process(R_MAX_COUNT_9434_wire_constant, count_9432) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(R_MAX_COUNT_9434_wire_constant, count_9432, tmp_var);
      ULT_u15_u1_9436_wire <= tmp_var; -- 
    end process;
    -- binary operator ULT_u15_u1_9474_inst
    process(count_var_9449, count_blocks_9447) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(count_var_9449, count_blocks_9447, tmp_var);
      ULT_u15_u1_9474_wire <= tmp_var; -- 
    end process;
    -- binary operator ULT_u15_u1_9480_inst
    process(count_var_9449) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(count_var_9449, R_MAX_COUNT_9479_wire_constant, tmp_var);
      ULT_u15_u1_9480_wire <= tmp_var; -- 
    end process;
    -- binary operator ULT_u15_u1_9498_inst
    process(count_var2_9482) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(count_var2_9482, R_MAX_COUNT_9497_wire_constant, tmp_var);
      ULT_u15_u1_9498_wire <= tmp_var; -- 
    end process;
    -- shared inport operator group (0) : RPIPE_d_out_buf_9463_inst 
    InportGroup0: Block -- 
      signal data_out: std_logic_vector(127 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_d_out_buf_9463_inst_req_0;
      RPIPE_d_out_buf_9463_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_d_out_buf_9463_inst_req_1;
      RPIPE_d_out_buf_9463_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      gI: SplitGuardInterface generic map(name => "gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      RPIPE_d_out_buf_9463_wire <= data_out(127 downto 0);
      d_out_buf_read_0: InputPortRevised -- 
        generic map ( name => "d_out_buf_read_0", data_width => 128,  num_reqs => 1,  output_buffering => outBUFs,   no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => d_out_buf_pipe_read_req(0),
          oack => d_out_buf_pipe_read_ack(0),
          odata => d_out_buf_pipe_read_data(127 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared inport operator group (1) : RPIPE_e_out_buf_9459_inst 
    InportGroup1: Block -- 
      signal data_out: std_logic_vector(127 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_e_out_buf_9459_inst_req_0;
      RPIPE_e_out_buf_9459_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_e_out_buf_9459_inst_req_1;
      RPIPE_e_out_buf_9459_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      gI: SplitGuardInterface generic map(name => "gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      RPIPE_e_out_buf_9459_wire <= data_out(127 downto 0);
      e_out_buf_read_1: InputPortRevised -- 
        generic map ( name => "e_out_buf_read_1", data_width => 128,  num_reqs => 1,  output_buffering => outBUFs,   no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => e_out_buf_pipe_read_req(0),
          oack => e_out_buf_pipe_read_ack(0),
          odata => e_out_buf_pipe_read_data(127 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 1
    -- shared inport operator group (2) : RPIPE_out_wrap_cmd_9403_inst 
    InportGroup2: Block -- 
      signal data_out: std_logic_vector(63 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_out_wrap_cmd_9403_inst_req_0;
      RPIPE_out_wrap_cmd_9403_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_out_wrap_cmd_9403_inst_req_1;
      RPIPE_out_wrap_cmd_9403_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      gI: SplitGuardInterface generic map(name => "gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      head_out_9404 <= data_out(63 downto 0);
      out_wrap_cmd_read_2: InputPortRevised -- 
        generic map ( name => "out_wrap_cmd_read_2", data_width => 64,  num_reqs => 1,  output_buffering => outBUFs,   no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => out_wrap_cmd_pipe_read_req(0),
          oack => out_wrap_cmd_pipe_read_ack(0),
          odata => out_wrap_cmd_pipe_read_data(63 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 2
    -- shared inport operator group (3) : RPIPE_out_wrap_data_9488_inst 
    InportGroup3: Block -- 
      signal data_out: std_logic_vector(127 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_out_wrap_data_9488_inst_req_0;
      RPIPE_out_wrap_data_9488_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_out_wrap_data_9488_inst_req_1;
      RPIPE_out_wrap_data_9488_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      gI: SplitGuardInterface generic map(name => "gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      RPIPE_out_wrap_data_9488_wire <= data_out(127 downto 0);
      out_wrap_data_read_3: InputPortRevised -- 
        generic map ( name => "out_wrap_data_read_3", data_width => 128,  num_reqs => 1,  output_buffering => outBUFs,   no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => out_wrap_data_pipe_read_req(0),
          oack => out_wrap_data_pipe_read_ack(0),
          odata => out_wrap_data_pipe_read_data(127 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 3
    -- shared inport operator group (4) : RPIPE_status_out_9406_inst 
    InportGroup4: Block -- 
      signal data_out: std_logic_vector(63 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_status_out_9406_inst_req_0;
      RPIPE_status_out_9406_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_status_out_9406_inst_req_1;
      RPIPE_status_out_9406_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      gI: SplitGuardInterface generic map(name => "gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      st_out_9407 <= data_out(63 downto 0);
      status_out_read_4: InputPortRevised -- 
        generic map ( name => "status_out_read_4", data_width => 64,  num_reqs => 1,  output_buffering => outBUFs,   no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => status_out_pipe_read_req(0),
          oack => status_out_pipe_read_ack(0),
          odata => status_out_pipe_read_data(63 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 4
    -- shared outport operator group (0) : WPIPE_w_out_buf_9408_inst WPIPE_w_out_buf_9462_inst WPIPE_w_out_buf_9458_inst WPIPE_w_out_buf_9487_inst 
    OutportGroup0: Block -- 
      signal data_in: std_logic_vector(511 downto 0);
      signal sample_req, sample_ack : BooleanArray( 3 downto 0);
      signal update_req, update_ack : BooleanArray( 3 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 3 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 3 downto 0);
      signal guard_vector : std_logic_vector( 3 downto 0);
      constant inBUFs : IntegerArray(3 downto 0) := (3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(3 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false);
      constant guardBuffering: IntegerArray(3 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2);
      -- 
    begin -- 
      sample_req_unguarded(3) <= WPIPE_w_out_buf_9408_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_w_out_buf_9462_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_w_out_buf_9458_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_w_out_buf_9487_inst_req_0;
      WPIPE_w_out_buf_9408_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_w_out_buf_9462_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_w_out_buf_9458_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_w_out_buf_9487_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(3) <= WPIPE_w_out_buf_9408_inst_req_1;
      update_req_unguarded(2) <= WPIPE_w_out_buf_9462_inst_req_1;
      update_req_unguarded(1) <= WPIPE_w_out_buf_9458_inst_req_1;
      update_req_unguarded(0) <= WPIPE_w_out_buf_9487_inst_req_1;
      WPIPE_w_out_buf_9408_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_w_out_buf_9462_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_w_out_buf_9458_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_w_out_buf_9487_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      gI: SplitGuardInterface generic map(name => "gI", nreqs => 4, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      data_in <= CONCAT_u64_u128_9411_wire & RPIPE_d_out_buf_9463_wire & RPIPE_e_out_buf_9459_wire & RPIPE_out_wrap_data_9488_wire;
      w_out_buf_write_0: OutputPortRevised -- 
        generic map ( name => "w_out_buf", data_width => 128, num_reqs => 4, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => w_out_buf_pipe_write_req(0),
          oack => w_out_buf_pipe_write_ack(0),
          odata => w_out_buf_pipe_write_data(127 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end Out_wrap_daemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library work;
use work.ahir_system_global_package.all;
entity c_block_daemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    cmd_in_pipe_read_req : out  std_logic_vector(0 downto 0);
    cmd_in_pipe_read_ack : in   std_logic_vector(0 downto 0);
    cmd_in_pipe_read_data : in   std_logic_vector(63 downto 0);
    d_block_done_pipe_read_req : out  std_logic_vector(0 downto 0);
    d_block_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
    d_block_done_pipe_read_data : in   std_logic_vector(0 downto 0);
    e_block_done_pipe_read_req : out  std_logic_vector(0 downto 0);
    e_block_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
    e_block_done_pipe_read_data : in   std_logic_vector(0 downto 0);
    d_cmd_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    d_cmd_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    d_cmd_pipe_pipe_write_data : out  std_logic_vector(143 downto 0);
    e_cmd_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    e_cmd_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    e_cmd_pipe_pipe_write_data : out  std_logic_vector(143 downto 0);
    status_out_pipe_write_req : out  std_logic_vector(0 downto 0);
    status_out_pipe_write_ack : in   std_logic_vector(0 downto 0);
    status_out_pipe_write_data : out  std_logic_vector(63 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity c_block_daemon;
architecture c_block_daemon_arch of c_block_daemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal c_block_daemon_CP_1519_start: Boolean;
  signal c_block_daemon_CP_1519_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal RPIPE_d_block_done_9579_inst_req_1 : boolean;
  signal RPIPE_d_block_done_9579_inst_ack_1 : boolean;
  signal if_stmt_9581_branch_ack_0 : boolean;
  signal if_stmt_9581_branch_ack_1 : boolean;
  signal if_stmt_9581_branch_req_0 : boolean;
  signal WPIPE_status_out_9574_inst_ack_1 : boolean;
  signal RPIPE_d_block_done_9579_inst_ack_0 : boolean;
  signal if_stmt_9570_branch_ack_0 : boolean;
  signal if_stmt_9570_branch_ack_1 : boolean;
  signal RPIPE_d_block_done_9579_inst_req_0 : boolean;
  signal WPIPE_status_out_9574_inst_req_1 : boolean;
  signal WPIPE_status_out_9574_inst_ack_0 : boolean;
  signal WPIPE_status_out_9574_inst_req_0 : boolean;
  signal if_stmt_9570_branch_req_0 : boolean;
  signal RPIPE_cmd_in_9507_inst_req_0 : boolean;
  signal RPIPE_cmd_in_9507_inst_ack_0 : boolean;
  signal RPIPE_cmd_in_9507_inst_req_1 : boolean;
  signal RPIPE_cmd_in_9507_inst_ack_1 : boolean;
  signal RPIPE_cmd_in_9530_inst_req_0 : boolean;
  signal RPIPE_cmd_in_9530_inst_ack_0 : boolean;
  signal RPIPE_cmd_in_9530_inst_req_1 : boolean;
  signal RPIPE_cmd_in_9530_inst_ack_1 : boolean;
  signal RPIPE_cmd_in_9534_inst_req_0 : boolean;
  signal RPIPE_cmd_in_9534_inst_ack_0 : boolean;
  signal RPIPE_cmd_in_9534_inst_req_1 : boolean;
  signal RPIPE_cmd_in_9534_inst_ack_1 : boolean;
  signal if_stmt_9538_branch_req_0 : boolean;
  signal if_stmt_9538_branch_ack_1 : boolean;
  signal if_stmt_9538_branch_ack_0 : boolean;
  signal WPIPE_status_out_9542_inst_req_0 : boolean;
  signal WPIPE_status_out_9542_inst_ack_0 : boolean;
  signal WPIPE_status_out_9542_inst_req_1 : boolean;
  signal WPIPE_status_out_9542_inst_ack_1 : boolean;
  signal RPIPE_e_block_done_9547_inst_req_0 : boolean;
  signal RPIPE_e_block_done_9547_inst_ack_0 : boolean;
  signal RPIPE_e_block_done_9547_inst_req_1 : boolean;
  signal RPIPE_e_block_done_9547_inst_ack_1 : boolean;
  signal if_stmt_9549_branch_req_0 : boolean;
  signal if_stmt_9549_branch_ack_1 : boolean;
  signal if_stmt_9549_branch_ack_0 : boolean;
  signal WPIPE_e_cmd_pipe_9564_inst_req_0 : boolean;
  signal WPIPE_e_cmd_pipe_9564_inst_ack_0 : boolean;
  signal WPIPE_e_cmd_pipe_9564_inst_req_1 : boolean;
  signal WPIPE_e_cmd_pipe_9564_inst_ack_1 : boolean;
  signal WPIPE_d_cmd_pipe_9596_inst_req_0 : boolean;
  signal WPIPE_d_cmd_pipe_9596_inst_ack_0 : boolean;
  signal WPIPE_d_cmd_pipe_9596_inst_req_1 : boolean;
  signal WPIPE_d_cmd_pipe_9596_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "c_block_daemon_input_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      bypass_flag => true,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  c_block_daemon_CP_1519_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "c_block_daemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= c_block_daemon_CP_1519_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= c_block_daemon_CP_1519_start & tag_ilock_write_ack_symbol;
    gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= c_block_daemon_CP_1519_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  c_block_daemon_CP_1519: Block -- control-path 
    signal c_block_daemon_CP_1519_elements: BooleanArray(88 downto 0);
    -- 
  begin -- 
    c_block_daemon_CP_1519_elements(0) <= c_block_daemon_CP_1519_start;
    c_block_daemon_CP_1519_symbol <= c_block_daemon_CP_1519_elements(88);
    -- CP-element group 0:  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (5) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_9508/$entry
      -- CP-element group 0: 	 assign_stmt_9508/RPIPE_cmd_in_9507_sample_start_
      -- CP-element group 0: 	 assign_stmt_9508/RPIPE_cmd_in_9507_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_9508/RPIPE_cmd_in_9507_Sample/rr
      -- 
    rr_1532_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1532_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => c_block_daemon_CP_1519_elements(0), ack => RPIPE_cmd_in_9507_inst_req_0); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 assign_stmt_9508/RPIPE_cmd_in_9507_sample_completed_
      -- CP-element group 1: 	 assign_stmt_9508/RPIPE_cmd_in_9507_update_start_
      -- CP-element group 1: 	 assign_stmt_9508/RPIPE_cmd_in_9507_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_9508/RPIPE_cmd_in_9507_Sample/ra
      -- CP-element group 1: 	 assign_stmt_9508/RPIPE_cmd_in_9507_Update/$entry
      -- CP-element group 1: 	 assign_stmt_9508/RPIPE_cmd_in_9507_Update/cr
      -- 
    ra_1533_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_cmd_in_9507_inst_ack_0, ack => c_block_daemon_CP_1519_elements(1)); -- 
    cr_1537_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1537_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => c_block_daemon_CP_1519_elements(1), ack => RPIPE_cmd_in_9507_inst_req_1); -- 
    -- CP-element group 2:  join  fork  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2: 	5 
    -- CP-element group 2:  members (94) 
      -- CP-element group 2: 	 assign_stmt_9508/$exit
      -- CP-element group 2: 	 assign_stmt_9508/RPIPE_cmd_in_9507_update_completed_
      -- CP-element group 2: 	 assign_stmt_9508/RPIPE_cmd_in_9507_Update/$exit
      -- CP-element group 2: 	 assign_stmt_9508/RPIPE_cmd_in_9507_Update/ca
      -- CP-element group 2: 	 assign_stmt_9512_to_assign_stmt_9528/$entry
      -- CP-element group 2: 	 assign_stmt_9512_to_assign_stmt_9528/$exit
      -- CP-element group 2: 	 assign_stmt_9512_to_assign_stmt_9528/slice_9511_sample_start_
      -- CP-element group 2: 	 assign_stmt_9512_to_assign_stmt_9528/slice_9511_sample_completed_
      -- CP-element group 2: 	 assign_stmt_9512_to_assign_stmt_9528/slice_9511_update_start_
      -- CP-element group 2: 	 assign_stmt_9512_to_assign_stmt_9528/slice_9511_update_completed_
      -- CP-element group 2: 	 assign_stmt_9512_to_assign_stmt_9528/R_command_9510_sample_start_
      -- CP-element group 2: 	 assign_stmt_9512_to_assign_stmt_9528/R_command_9510_sample_completed_
      -- CP-element group 2: 	 assign_stmt_9512_to_assign_stmt_9528/R_command_9510_update_start_
      -- CP-element group 2: 	 assign_stmt_9512_to_assign_stmt_9528/R_command_9510_update_completed_
      -- CP-element group 2: 	 assign_stmt_9512_to_assign_stmt_9528/slice_9511_Sample/$entry
      -- CP-element group 2: 	 assign_stmt_9512_to_assign_stmt_9528/slice_9511_Sample/$exit
      -- CP-element group 2: 	 assign_stmt_9512_to_assign_stmt_9528/slice_9511_Sample/rr
      -- CP-element group 2: 	 assign_stmt_9512_to_assign_stmt_9528/slice_9511_Sample/ra
      -- CP-element group 2: 	 assign_stmt_9512_to_assign_stmt_9528/slice_9511_Update/$entry
      -- CP-element group 2: 	 assign_stmt_9512_to_assign_stmt_9528/slice_9511_Update/$exit
      -- CP-element group 2: 	 assign_stmt_9512_to_assign_stmt_9528/slice_9511_Update/cr
      -- CP-element group 2: 	 assign_stmt_9512_to_assign_stmt_9528/slice_9511_Update/ca
      -- CP-element group 2: 	 assign_stmt_9512_to_assign_stmt_9528/slice_9515_sample_start_
      -- CP-element group 2: 	 assign_stmt_9512_to_assign_stmt_9528/slice_9515_sample_completed_
      -- CP-element group 2: 	 assign_stmt_9512_to_assign_stmt_9528/slice_9515_update_start_
      -- CP-element group 2: 	 assign_stmt_9512_to_assign_stmt_9528/slice_9515_update_completed_
      -- CP-element group 2: 	 assign_stmt_9512_to_assign_stmt_9528/R_command_9514_sample_start_
      -- CP-element group 2: 	 assign_stmt_9512_to_assign_stmt_9528/R_command_9514_sample_completed_
      -- CP-element group 2: 	 assign_stmt_9512_to_assign_stmt_9528/R_command_9514_update_start_
      -- CP-element group 2: 	 assign_stmt_9512_to_assign_stmt_9528/R_command_9514_update_completed_
      -- CP-element group 2: 	 assign_stmt_9512_to_assign_stmt_9528/slice_9515_Sample/$entry
      -- CP-element group 2: 	 assign_stmt_9512_to_assign_stmt_9528/slice_9515_Sample/$exit
      -- CP-element group 2: 	 assign_stmt_9512_to_assign_stmt_9528/slice_9515_Sample/rr
      -- CP-element group 2: 	 assign_stmt_9512_to_assign_stmt_9528/slice_9515_Sample/ra
      -- CP-element group 2: 	 assign_stmt_9512_to_assign_stmt_9528/slice_9515_Update/$entry
      -- CP-element group 2: 	 assign_stmt_9512_to_assign_stmt_9528/slice_9515_Update/$exit
      -- CP-element group 2: 	 assign_stmt_9512_to_assign_stmt_9528/slice_9515_Update/cr
      -- CP-element group 2: 	 assign_stmt_9512_to_assign_stmt_9528/slice_9515_Update/ca
      -- CP-element group 2: 	 assign_stmt_9512_to_assign_stmt_9528/slice_9519_sample_start_
      -- CP-element group 2: 	 assign_stmt_9512_to_assign_stmt_9528/slice_9519_sample_completed_
      -- CP-element group 2: 	 assign_stmt_9512_to_assign_stmt_9528/slice_9519_update_start_
      -- CP-element group 2: 	 assign_stmt_9512_to_assign_stmt_9528/slice_9519_update_completed_
      -- CP-element group 2: 	 assign_stmt_9512_to_assign_stmt_9528/R_command_9518_sample_start_
      -- CP-element group 2: 	 assign_stmt_9512_to_assign_stmt_9528/R_command_9518_sample_completed_
      -- CP-element group 2: 	 assign_stmt_9512_to_assign_stmt_9528/R_command_9518_update_start_
      -- CP-element group 2: 	 assign_stmt_9512_to_assign_stmt_9528/R_command_9518_update_completed_
      -- CP-element group 2: 	 assign_stmt_9512_to_assign_stmt_9528/slice_9519_Sample/$entry
      -- CP-element group 2: 	 assign_stmt_9512_to_assign_stmt_9528/slice_9519_Sample/$exit
      -- CP-element group 2: 	 assign_stmt_9512_to_assign_stmt_9528/slice_9519_Sample/rr
      -- CP-element group 2: 	 assign_stmt_9512_to_assign_stmt_9528/slice_9519_Sample/ra
      -- CP-element group 2: 	 assign_stmt_9512_to_assign_stmt_9528/slice_9519_Update/$entry
      -- CP-element group 2: 	 assign_stmt_9512_to_assign_stmt_9528/slice_9519_Update/$exit
      -- CP-element group 2: 	 assign_stmt_9512_to_assign_stmt_9528/slice_9519_Update/cr
      -- CP-element group 2: 	 assign_stmt_9512_to_assign_stmt_9528/slice_9519_Update/ca
      -- CP-element group 2: 	 assign_stmt_9512_to_assign_stmt_9528/slice_9523_sample_start_
      -- CP-element group 2: 	 assign_stmt_9512_to_assign_stmt_9528/slice_9523_sample_completed_
      -- CP-element group 2: 	 assign_stmt_9512_to_assign_stmt_9528/slice_9523_update_start_
      -- CP-element group 2: 	 assign_stmt_9512_to_assign_stmt_9528/slice_9523_update_completed_
      -- CP-element group 2: 	 assign_stmt_9512_to_assign_stmt_9528/R_command_9522_sample_start_
      -- CP-element group 2: 	 assign_stmt_9512_to_assign_stmt_9528/R_command_9522_sample_completed_
      -- CP-element group 2: 	 assign_stmt_9512_to_assign_stmt_9528/R_command_9522_update_start_
      -- CP-element group 2: 	 assign_stmt_9512_to_assign_stmt_9528/R_command_9522_update_completed_
      -- CP-element group 2: 	 assign_stmt_9512_to_assign_stmt_9528/slice_9523_Sample/$entry
      -- CP-element group 2: 	 assign_stmt_9512_to_assign_stmt_9528/slice_9523_Sample/$exit
      -- CP-element group 2: 	 assign_stmt_9512_to_assign_stmt_9528/slice_9523_Sample/rr
      -- CP-element group 2: 	 assign_stmt_9512_to_assign_stmt_9528/slice_9523_Sample/ra
      -- CP-element group 2: 	 assign_stmt_9512_to_assign_stmt_9528/slice_9523_Update/$entry
      -- CP-element group 2: 	 assign_stmt_9512_to_assign_stmt_9528/slice_9523_Update/$exit
      -- CP-element group 2: 	 assign_stmt_9512_to_assign_stmt_9528/slice_9523_Update/cr
      -- CP-element group 2: 	 assign_stmt_9512_to_assign_stmt_9528/slice_9523_Update/ca
      -- CP-element group 2: 	 assign_stmt_9512_to_assign_stmt_9528/slice_9527_sample_start_
      -- CP-element group 2: 	 assign_stmt_9512_to_assign_stmt_9528/slice_9527_sample_completed_
      -- CP-element group 2: 	 assign_stmt_9512_to_assign_stmt_9528/slice_9527_update_start_
      -- CP-element group 2: 	 assign_stmt_9512_to_assign_stmt_9528/slice_9527_update_completed_
      -- CP-element group 2: 	 assign_stmt_9512_to_assign_stmt_9528/R_command_9526_sample_start_
      -- CP-element group 2: 	 assign_stmt_9512_to_assign_stmt_9528/R_command_9526_sample_completed_
      -- CP-element group 2: 	 assign_stmt_9512_to_assign_stmt_9528/R_command_9526_update_start_
      -- CP-element group 2: 	 assign_stmt_9512_to_assign_stmt_9528/R_command_9526_update_completed_
      -- CP-element group 2: 	 assign_stmt_9512_to_assign_stmt_9528/slice_9527_Sample/$entry
      -- CP-element group 2: 	 assign_stmt_9512_to_assign_stmt_9528/slice_9527_Sample/$exit
      -- CP-element group 2: 	 assign_stmt_9512_to_assign_stmt_9528/slice_9527_Sample/rr
      -- CP-element group 2: 	 assign_stmt_9512_to_assign_stmt_9528/slice_9527_Sample/ra
      -- CP-element group 2: 	 assign_stmt_9512_to_assign_stmt_9528/slice_9527_Update/$entry
      -- CP-element group 2: 	 assign_stmt_9512_to_assign_stmt_9528/slice_9527_Update/$exit
      -- CP-element group 2: 	 assign_stmt_9512_to_assign_stmt_9528/slice_9527_Update/cr
      -- CP-element group 2: 	 assign_stmt_9512_to_assign_stmt_9528/slice_9527_Update/ca
      -- CP-element group 2: 	 assign_stmt_9531/$entry
      -- CP-element group 2: 	 assign_stmt_9531/R_got_new_key_9532_sample_start_
      -- CP-element group 2: 	 assign_stmt_9531/R_got_new_key_9532_sample_completed_
      -- CP-element group 2: 	 assign_stmt_9531/R_got_new_key_9532_update_start_
      -- CP-element group 2: 	 assign_stmt_9531/R_got_new_key_9532_update_completed_
      -- CP-element group 2: 	 assign_stmt_9531/RPIPE_cmd_in_9530_sample_start_
      -- CP-element group 2: 	 assign_stmt_9531/RPIPE_cmd_in_9530_Sample/$entry
      -- CP-element group 2: 	 assign_stmt_9531/RPIPE_cmd_in_9530_Sample/rr
      -- 
    ca_1538_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_cmd_in_9507_inst_ack_1, ack => c_block_daemon_CP_1519_elements(2)); -- 
    rr_1646_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1646_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => c_block_daemon_CP_1519_elements(2), ack => RPIPE_cmd_in_9530_inst_req_0); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 assign_stmt_9531/RPIPE_cmd_in_9530_sample_completed_
      -- CP-element group 3: 	 assign_stmt_9531/RPIPE_cmd_in_9530_update_start_
      -- CP-element group 3: 	 assign_stmt_9531/RPIPE_cmd_in_9530_Sample/$exit
      -- CP-element group 3: 	 assign_stmt_9531/RPIPE_cmd_in_9530_Sample/ra
      -- CP-element group 3: 	 assign_stmt_9531/RPIPE_cmd_in_9530_Update/$entry
      -- CP-element group 3: 	 assign_stmt_9531/RPIPE_cmd_in_9530_Update/cr
      -- 
    ra_1647_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_cmd_in_9530_inst_ack_0, ack => c_block_daemon_CP_1519_elements(3)); -- 
    cr_1651_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1651_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => c_block_daemon_CP_1519_elements(3), ack => RPIPE_cmd_in_9530_inst_req_1); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 assign_stmt_9531/RPIPE_cmd_in_9530_update_completed_
      -- CP-element group 4: 	 assign_stmt_9531/RPIPE_cmd_in_9530_Update/$exit
      -- CP-element group 4: 	 assign_stmt_9531/RPIPE_cmd_in_9530_Update/ca
      -- 
    ca_1652_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_cmd_in_9530_inst_ack_1, ack => c_block_daemon_CP_1519_elements(4)); -- 
    -- CP-element group 5:  join  fork  transition  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	2 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5: 	8 
    -- CP-element group 5:  members (9) 
      -- CP-element group 5: 	 assign_stmt_9531/$exit
      -- CP-element group 5: 	 assign_stmt_9535/$entry
      -- CP-element group 5: 	 assign_stmt_9535/R_got_new_key_9536_sample_start_
      -- CP-element group 5: 	 assign_stmt_9535/R_got_new_key_9536_sample_completed_
      -- CP-element group 5: 	 assign_stmt_9535/R_got_new_key_9536_update_start_
      -- CP-element group 5: 	 assign_stmt_9535/R_got_new_key_9536_update_completed_
      -- CP-element group 5: 	 assign_stmt_9535/RPIPE_cmd_in_9534_sample_start_
      -- CP-element group 5: 	 assign_stmt_9535/RPIPE_cmd_in_9534_Sample/$entry
      -- CP-element group 5: 	 assign_stmt_9535/RPIPE_cmd_in_9534_Sample/rr
      -- 
    rr_1667_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1667_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => c_block_daemon_CP_1519_elements(5), ack => RPIPE_cmd_in_9534_inst_req_0); -- 
    c_block_daemon_cp_element_group_5: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "c_block_daemon_cp_element_group_5"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= c_block_daemon_CP_1519_elements(2) & c_block_daemon_CP_1519_elements(4);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => c_block_daemon_CP_1519_elements(5), clk => clk, reset => reset); --
    end block;
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (6) 
      -- CP-element group 6: 	 assign_stmt_9535/RPIPE_cmd_in_9534_sample_completed_
      -- CP-element group 6: 	 assign_stmt_9535/RPIPE_cmd_in_9534_update_start_
      -- CP-element group 6: 	 assign_stmt_9535/RPIPE_cmd_in_9534_Sample/$exit
      -- CP-element group 6: 	 assign_stmt_9535/RPIPE_cmd_in_9534_Sample/ra
      -- CP-element group 6: 	 assign_stmt_9535/RPIPE_cmd_in_9534_Update/$entry
      -- CP-element group 6: 	 assign_stmt_9535/RPIPE_cmd_in_9534_Update/cr
      -- 
    ra_1668_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_cmd_in_9534_inst_ack_0, ack => c_block_daemon_CP_1519_elements(6)); -- 
    cr_1672_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1672_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => c_block_daemon_CP_1519_elements(6), ack => RPIPE_cmd_in_9534_inst_req_1); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 assign_stmt_9535/RPIPE_cmd_in_9534_update_completed_
      -- CP-element group 7: 	 assign_stmt_9535/RPIPE_cmd_in_9534_Update/$exit
      -- CP-element group 7: 	 assign_stmt_9535/RPIPE_cmd_in_9534_Update/ca
      -- 
    ca_1673_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_cmd_in_9534_inst_ack_1, ack => c_block_daemon_CP_1519_elements(7)); -- 
    -- CP-element group 8:  join  transition  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	5 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (2) 
      -- CP-element group 8: 	 assign_stmt_9535/$exit
      -- CP-element group 8: 	 branch_block_stmt_9537/$entry
      -- 
    c_block_daemon_cp_element_group_8: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "c_block_daemon_cp_element_group_8"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= c_block_daemon_CP_1519_elements(5) & c_block_daemon_CP_1519_elements(7);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => c_block_daemon_CP_1519_elements(8), clk => clk, reset => reset); --
    end block;
    -- CP-element group 9:  branch  place  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	11 
    -- CP-element group 9: 	12 
    -- CP-element group 9:  members (2) 
      -- CP-element group 9: 	 branch_block_stmt_9537/branch_block_stmt_9537__entry__
      -- CP-element group 9: 	 branch_block_stmt_9537/if_stmt_9538__entry__
      -- 
    c_block_daemon_CP_1519_elements(9) <= c_block_daemon_CP_1519_elements(8);
    -- CP-element group 10:  merge  place  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	17 
    -- CP-element group 10: 	24 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	48 
    -- CP-element group 10:  members (2) 
      -- CP-element group 10: 	 branch_block_stmt_9537/branch_block_stmt_9537__exit__
      -- CP-element group 10: 	 branch_block_stmt_9537/if_stmt_9538__exit__
      -- 
    c_block_daemon_CP_1519_elements(10) <= OrReduce(c_block_daemon_CP_1519_elements(17) & c_block_daemon_CP_1519_elements(24));
    -- CP-element group 11:  transition  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (1) 
      -- CP-element group 11: 	 branch_block_stmt_9537/if_stmt_9538_dead_link/$entry
      -- 
    c_block_daemon_CP_1519_elements(11) <= c_block_daemon_CP_1519_elements(9);
    -- CP-element group 12:  transition  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	9 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (17) 
      -- CP-element group 12: 	 branch_block_stmt_9537/if_stmt_9538_eval_test/$entry
      -- CP-element group 12: 	 branch_block_stmt_9537/if_stmt_9538_eval_test/$exit
      -- CP-element group 12: 	 branch_block_stmt_9537/if_stmt_9538_eval_test/EQ_u1_u1_9541/$entry
      -- CP-element group 12: 	 branch_block_stmt_9537/if_stmt_9538_eval_test/EQ_u1_u1_9541/$exit
      -- CP-element group 12: 	 branch_block_stmt_9537/if_stmt_9538_eval_test/EQ_u1_u1_9541/EQ_u1_u1_9541_inputs/$entry
      -- CP-element group 12: 	 branch_block_stmt_9537/if_stmt_9538_eval_test/EQ_u1_u1_9541/EQ_u1_u1_9541_inputs/$exit
      -- CP-element group 12: 	 branch_block_stmt_9537/if_stmt_9538_eval_test/EQ_u1_u1_9541/SplitProtocol/$entry
      -- CP-element group 12: 	 branch_block_stmt_9537/if_stmt_9538_eval_test/EQ_u1_u1_9541/SplitProtocol/$exit
      -- CP-element group 12: 	 branch_block_stmt_9537/if_stmt_9538_eval_test/EQ_u1_u1_9541/SplitProtocol/Sample/$entry
      -- CP-element group 12: 	 branch_block_stmt_9537/if_stmt_9538_eval_test/EQ_u1_u1_9541/SplitProtocol/Sample/$exit
      -- CP-element group 12: 	 branch_block_stmt_9537/if_stmt_9538_eval_test/EQ_u1_u1_9541/SplitProtocol/Sample/rr
      -- CP-element group 12: 	 branch_block_stmt_9537/if_stmt_9538_eval_test/EQ_u1_u1_9541/SplitProtocol/Sample/ra
      -- CP-element group 12: 	 branch_block_stmt_9537/if_stmt_9538_eval_test/EQ_u1_u1_9541/SplitProtocol/Update/$entry
      -- CP-element group 12: 	 branch_block_stmt_9537/if_stmt_9538_eval_test/EQ_u1_u1_9541/SplitProtocol/Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_9537/if_stmt_9538_eval_test/EQ_u1_u1_9541/SplitProtocol/Update/cr
      -- CP-element group 12: 	 branch_block_stmt_9537/if_stmt_9538_eval_test/EQ_u1_u1_9541/SplitProtocol/Update/ca
      -- CP-element group 12: 	 branch_block_stmt_9537/if_stmt_9538_eval_test/branch_req
      -- 
    branch_req_1707_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1707_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => c_block_daemon_CP_1519_elements(12), ack => if_stmt_9538_branch_req_0); -- 
    c_block_daemon_CP_1519_elements(12) <= c_block_daemon_CP_1519_elements(9);
    -- CP-element group 13:  branch  place  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13: 	16 
    -- CP-element group 13:  members (1) 
      -- CP-element group 13: 	 branch_block_stmt_9537/EQ_u1_u1_9541_place
      -- 
    c_block_daemon_CP_1519_elements(13) <= c_block_daemon_CP_1519_elements(12);
    -- CP-element group 14:  transition  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 branch_block_stmt_9537/if_stmt_9538_if_link/$entry
      -- 
    c_block_daemon_CP_1519_elements(14) <= c_block_daemon_CP_1519_elements(13);
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	18 
    -- CP-element group 15:  members (2) 
      -- CP-element group 15: 	 branch_block_stmt_9537/if_stmt_9538_if_link/$exit
      -- CP-element group 15: 	 branch_block_stmt_9537/if_stmt_9538_if_link/if_choice_transition
      -- 
    if_choice_transition_1712_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_9538_branch_ack_1, ack => c_block_daemon_CP_1519_elements(15)); -- 
    -- CP-element group 16:  transition  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	13 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	17 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_9537/if_stmt_9538_else_link/$entry
      -- 
    c_block_daemon_CP_1519_elements(16) <= c_block_daemon_CP_1519_elements(13);
    -- CP-element group 17:  transition  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	16 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	10 
    -- CP-element group 17:  members (2) 
      -- CP-element group 17: 	 branch_block_stmt_9537/if_stmt_9538_else_link/$exit
      -- CP-element group 17: 	 branch_block_stmt_9537/if_stmt_9538_else_link/else_choice_transition
      -- 
    else_choice_transition_1716_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_9538_branch_ack_0, ack => c_block_daemon_CP_1519_elements(17)); -- 
    -- CP-element group 18:  place  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	15 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	25 
    -- CP-element group 18:  members (1) 
      -- CP-element group 18: 	 branch_block_stmt_9537/assign_stmt_9544__entry__
      -- 
    c_block_daemon_CP_1519_elements(18) <= c_block_daemon_CP_1519_elements(15);
    -- CP-element group 19:  branch  place  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	27 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	43 
    -- CP-element group 19: 	44 
    -- CP-element group 19:  members (2) 
      -- CP-element group 19: 	 branch_block_stmt_9537/assign_stmt_9544__exit__
      -- CP-element group 19: 	 branch_block_stmt_9537/merge_stmt_9545__entry__
      -- 
    c_block_daemon_CP_1519_elements(19) <= c_block_daemon_CP_1519_elements(27);
    -- CP-element group 20:  merge  place  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	47 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	28 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_9537/merge_stmt_9545__exit__
      -- CP-element group 20: 	 branch_block_stmt_9537/assign_stmt_9548__entry__
      -- 
    c_block_daemon_CP_1519_elements(20) <= c_block_daemon_CP_1519_elements(47);
    -- CP-element group 21:  branch  place  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	30 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	31 
    -- CP-element group 21: 	32 
    -- CP-element group 21:  members (2) 
      -- CP-element group 21: 	 branch_block_stmt_9537/assign_stmt_9548__exit__
      -- CP-element group 21: 	 branch_block_stmt_9537/if_stmt_9549__entry__
      -- 
    c_block_daemon_CP_1519_elements(21) <= c_block_daemon_CP_1519_elements(30);
    -- CP-element group 22:  merge  place  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	37 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	39 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_9537/if_stmt_9549__exit__
      -- CP-element group 22: 	 branch_block_stmt_9537/assign_stmt_9563__entry__
      -- 
    c_block_daemon_CP_1519_elements(22) <= c_block_daemon_CP_1519_elements(37);
    -- CP-element group 23:  place  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	39 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	40 
    -- CP-element group 23:  members (2) 
      -- CP-element group 23: 	 branch_block_stmt_9537/assign_stmt_9563__exit__
      -- CP-element group 23: 	 branch_block_stmt_9537/assign_stmt_9566__entry__
      -- 
    c_block_daemon_CP_1519_elements(23) <= c_block_daemon_CP_1519_elements(39);
    -- CP-element group 24:  place  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	42 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	10 
    -- CP-element group 24:  members (1) 
      -- CP-element group 24: 	 branch_block_stmt_9537/assign_stmt_9566__exit__
      -- 
    c_block_daemon_CP_1519_elements(24) <= c_block_daemon_CP_1519_elements(42);
    -- CP-element group 25:  transition  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	18 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25:  members (4) 
      -- CP-element group 25: 	 branch_block_stmt_9537/assign_stmt_9544/$entry
      -- CP-element group 25: 	 branch_block_stmt_9537/assign_stmt_9544/WPIPE_status_out_9542_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_9537/assign_stmt_9544/WPIPE_status_out_9542_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_9537/assign_stmt_9544/WPIPE_status_out_9542_Sample/req
      -- 
    req_1739_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1739_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => c_block_daemon_CP_1519_elements(25), ack => WPIPE_status_out_9542_inst_req_0); -- 
    c_block_daemon_CP_1519_elements(25) <= c_block_daemon_CP_1519_elements(18);
    -- CP-element group 26:  transition  input  output  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	25 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	27 
    -- CP-element group 26:  members (6) 
      -- CP-element group 26: 	 branch_block_stmt_9537/assign_stmt_9544/WPIPE_status_out_9542_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_9537/assign_stmt_9544/WPIPE_status_out_9542_update_start_
      -- CP-element group 26: 	 branch_block_stmt_9537/assign_stmt_9544/WPIPE_status_out_9542_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_9537/assign_stmt_9544/WPIPE_status_out_9542_Sample/ack
      -- CP-element group 26: 	 branch_block_stmt_9537/assign_stmt_9544/WPIPE_status_out_9542_Update/$entry
      -- CP-element group 26: 	 branch_block_stmt_9537/assign_stmt_9544/WPIPE_status_out_9542_Update/req
      -- 
    ack_1740_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_status_out_9542_inst_ack_0, ack => c_block_daemon_CP_1519_elements(26)); -- 
    req_1744_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1744_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => c_block_daemon_CP_1519_elements(26), ack => WPIPE_status_out_9542_inst_req_1); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	26 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	19 
    -- CP-element group 27:  members (4) 
      -- CP-element group 27: 	 branch_block_stmt_9537/assign_stmt_9544/$exit
      -- CP-element group 27: 	 branch_block_stmt_9537/assign_stmt_9544/WPIPE_status_out_9542_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_9537/assign_stmt_9544/WPIPE_status_out_9542_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_9537/assign_stmt_9544/WPIPE_status_out_9542_Update/ack
      -- 
    ack_1745_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_status_out_9542_inst_ack_1, ack => c_block_daemon_CP_1519_elements(27)); -- 
    -- CP-element group 28:  transition  output  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	20 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28:  members (4) 
      -- CP-element group 28: 	 branch_block_stmt_9537/assign_stmt_9548/$entry
      -- CP-element group 28: 	 branch_block_stmt_9537/assign_stmt_9548/RPIPE_e_block_done_9547_sample_start_
      -- CP-element group 28: 	 branch_block_stmt_9537/assign_stmt_9548/RPIPE_e_block_done_9547_Sample/$entry
      -- CP-element group 28: 	 branch_block_stmt_9537/assign_stmt_9548/RPIPE_e_block_done_9547_Sample/rr
      -- 
    rr_1756_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1756_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => c_block_daemon_CP_1519_elements(28), ack => RPIPE_e_block_done_9547_inst_req_0); -- 
    c_block_daemon_CP_1519_elements(28) <= c_block_daemon_CP_1519_elements(20);
    -- CP-element group 29:  transition  input  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	28 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (6) 
      -- CP-element group 29: 	 branch_block_stmt_9537/assign_stmt_9548/RPIPE_e_block_done_9547_sample_completed_
      -- CP-element group 29: 	 branch_block_stmt_9537/assign_stmt_9548/RPIPE_e_block_done_9547_update_start_
      -- CP-element group 29: 	 branch_block_stmt_9537/assign_stmt_9548/RPIPE_e_block_done_9547_Sample/$exit
      -- CP-element group 29: 	 branch_block_stmt_9537/assign_stmt_9548/RPIPE_e_block_done_9547_Sample/ra
      -- CP-element group 29: 	 branch_block_stmt_9537/assign_stmt_9548/RPIPE_e_block_done_9547_Update/$entry
      -- CP-element group 29: 	 branch_block_stmt_9537/assign_stmt_9548/RPIPE_e_block_done_9547_Update/cr
      -- 
    ra_1757_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_e_block_done_9547_inst_ack_0, ack => c_block_daemon_CP_1519_elements(29)); -- 
    cr_1761_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1761_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => c_block_daemon_CP_1519_elements(29), ack => RPIPE_e_block_done_9547_inst_req_1); -- 
    -- CP-element group 30:  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	21 
    -- CP-element group 30:  members (4) 
      -- CP-element group 30: 	 branch_block_stmt_9537/assign_stmt_9548/$exit
      -- CP-element group 30: 	 branch_block_stmt_9537/assign_stmt_9548/RPIPE_e_block_done_9547_update_completed_
      -- CP-element group 30: 	 branch_block_stmt_9537/assign_stmt_9548/RPIPE_e_block_done_9547_Update/$exit
      -- CP-element group 30: 	 branch_block_stmt_9537/assign_stmt_9548/RPIPE_e_block_done_9547_Update/ca
      -- 
    ca_1762_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_e_block_done_9547_inst_ack_1, ack => c_block_daemon_CP_1519_elements(30)); -- 
    -- CP-element group 31:  transition  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	21 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (1) 
      -- CP-element group 31: 	 branch_block_stmt_9537/if_stmt_9549_dead_link/$entry
      -- 
    c_block_daemon_CP_1519_elements(31) <= c_block_daemon_CP_1519_elements(21);
    -- CP-element group 32:  transition  output  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	21 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	33 
    -- CP-element group 32:  members (17) 
      -- CP-element group 32: 	 branch_block_stmt_9537/if_stmt_9549_eval_test/$entry
      -- CP-element group 32: 	 branch_block_stmt_9537/if_stmt_9549_eval_test/$exit
      -- CP-element group 32: 	 branch_block_stmt_9537/if_stmt_9549_eval_test/EQ_u1_u1_9552/$entry
      -- CP-element group 32: 	 branch_block_stmt_9537/if_stmt_9549_eval_test/EQ_u1_u1_9552/$exit
      -- CP-element group 32: 	 branch_block_stmt_9537/if_stmt_9549_eval_test/EQ_u1_u1_9552/EQ_u1_u1_9552_inputs/$entry
      -- CP-element group 32: 	 branch_block_stmt_9537/if_stmt_9549_eval_test/EQ_u1_u1_9552/EQ_u1_u1_9552_inputs/$exit
      -- CP-element group 32: 	 branch_block_stmt_9537/if_stmt_9549_eval_test/EQ_u1_u1_9552/SplitProtocol/$entry
      -- CP-element group 32: 	 branch_block_stmt_9537/if_stmt_9549_eval_test/EQ_u1_u1_9552/SplitProtocol/$exit
      -- CP-element group 32: 	 branch_block_stmt_9537/if_stmt_9549_eval_test/EQ_u1_u1_9552/SplitProtocol/Sample/$entry
      -- CP-element group 32: 	 branch_block_stmt_9537/if_stmt_9549_eval_test/EQ_u1_u1_9552/SplitProtocol/Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_9537/if_stmt_9549_eval_test/EQ_u1_u1_9552/SplitProtocol/Sample/rr
      -- CP-element group 32: 	 branch_block_stmt_9537/if_stmt_9549_eval_test/EQ_u1_u1_9552/SplitProtocol/Sample/ra
      -- CP-element group 32: 	 branch_block_stmt_9537/if_stmt_9549_eval_test/EQ_u1_u1_9552/SplitProtocol/Update/$entry
      -- CP-element group 32: 	 branch_block_stmt_9537/if_stmt_9549_eval_test/EQ_u1_u1_9552/SplitProtocol/Update/$exit
      -- CP-element group 32: 	 branch_block_stmt_9537/if_stmt_9549_eval_test/EQ_u1_u1_9552/SplitProtocol/Update/cr
      -- CP-element group 32: 	 branch_block_stmt_9537/if_stmt_9549_eval_test/EQ_u1_u1_9552/SplitProtocol/Update/ca
      -- CP-element group 32: 	 branch_block_stmt_9537/if_stmt_9549_eval_test/branch_req
      -- 
    branch_req_1789_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1789_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => c_block_daemon_CP_1519_elements(32), ack => if_stmt_9549_branch_req_0); -- 
    c_block_daemon_CP_1519_elements(32) <= c_block_daemon_CP_1519_elements(21);
    -- CP-element group 33:  branch  place  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	32 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33: 	36 
    -- CP-element group 33:  members (1) 
      -- CP-element group 33: 	 branch_block_stmt_9537/EQ_u1_u1_9552_place
      -- 
    c_block_daemon_CP_1519_elements(33) <= c_block_daemon_CP_1519_elements(32);
    -- CP-element group 34:  transition  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34:  members (1) 
      -- CP-element group 34: 	 branch_block_stmt_9537/if_stmt_9549_if_link/$entry
      -- 
    c_block_daemon_CP_1519_elements(34) <= c_block_daemon_CP_1519_elements(33);
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	38 
    -- CP-element group 35:  members (2) 
      -- CP-element group 35: 	 branch_block_stmt_9537/if_stmt_9549_if_link/$exit
      -- CP-element group 35: 	 branch_block_stmt_9537/if_stmt_9549_if_link/if_choice_transition
      -- 
    if_choice_transition_1794_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_9549_branch_ack_1, ack => c_block_daemon_CP_1519_elements(35)); -- 
    -- CP-element group 36:  transition  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	33 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	37 
    -- CP-element group 36:  members (1) 
      -- CP-element group 36: 	 branch_block_stmt_9537/if_stmt_9549_else_link/$entry
      -- 
    c_block_daemon_CP_1519_elements(36) <= c_block_daemon_CP_1519_elements(33);
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	36 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	22 
    -- CP-element group 37:  members (2) 
      -- CP-element group 37: 	 branch_block_stmt_9537/if_stmt_9549_else_link/$exit
      -- CP-element group 37: 	 branch_block_stmt_9537/if_stmt_9549_else_link/else_choice_transition
      -- 
    else_choice_transition_1798_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_9549_branch_ack_0, ack => c_block_daemon_CP_1519_elements(37)); -- 
    -- CP-element group 38:  place  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	35 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	45 
    -- CP-element group 38:  members (1) 
      -- CP-element group 38: 	 branch_block_stmt_9537/e_block_BUSY
      -- 
    c_block_daemon_CP_1519_elements(38) <= c_block_daemon_CP_1519_elements(35);
    -- CP-element group 39:  join  fork  transition  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	22 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	23 
    -- CP-element group 39:  members (54) 
      -- CP-element group 39: 	 branch_block_stmt_9537/assign_stmt_9563/$entry
      -- CP-element group 39: 	 branch_block_stmt_9537/assign_stmt_9563/$exit
      -- CP-element group 39: 	 branch_block_stmt_9537/assign_stmt_9563/CONCAT_u16_u144_9562_sample_start_
      -- CP-element group 39: 	 branch_block_stmt_9537/assign_stmt_9563/CONCAT_u16_u144_9562_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_9537/assign_stmt_9563/CONCAT_u16_u144_9562_update_start_
      -- CP-element group 39: 	 branch_block_stmt_9537/assign_stmt_9563/CONCAT_u16_u144_9562_update_completed_
      -- CP-element group 39: 	 branch_block_stmt_9537/assign_stmt_9563/CONCAT_u1_u16_9558_sample_start_
      -- CP-element group 39: 	 branch_block_stmt_9537/assign_stmt_9563/CONCAT_u1_u16_9558_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_9537/assign_stmt_9563/CONCAT_u1_u16_9558_update_start_
      -- CP-element group 39: 	 branch_block_stmt_9537/assign_stmt_9563/CONCAT_u1_u16_9558_update_completed_
      -- CP-element group 39: 	 branch_block_stmt_9537/assign_stmt_9563/R_got_new_key_9556_sample_start_
      -- CP-element group 39: 	 branch_block_stmt_9537/assign_stmt_9563/R_got_new_key_9556_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_9537/assign_stmt_9563/R_got_new_key_9556_update_start_
      -- CP-element group 39: 	 branch_block_stmt_9537/assign_stmt_9563/R_got_new_key_9556_update_completed_
      -- CP-element group 39: 	 branch_block_stmt_9537/assign_stmt_9563/R_count_9557_sample_start_
      -- CP-element group 39: 	 branch_block_stmt_9537/assign_stmt_9563/R_count_9557_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_9537/assign_stmt_9563/R_count_9557_update_start_
      -- CP-element group 39: 	 branch_block_stmt_9537/assign_stmt_9563/R_count_9557_update_completed_
      -- CP-element group 39: 	 branch_block_stmt_9537/assign_stmt_9563/CONCAT_u1_u16_9558_Sample/$entry
      -- CP-element group 39: 	 branch_block_stmt_9537/assign_stmt_9563/CONCAT_u1_u16_9558_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_9537/assign_stmt_9563/CONCAT_u1_u16_9558_Sample/rr
      -- CP-element group 39: 	 branch_block_stmt_9537/assign_stmt_9563/CONCAT_u1_u16_9558_Sample/ra
      -- CP-element group 39: 	 branch_block_stmt_9537/assign_stmt_9563/CONCAT_u1_u16_9558_Update/$entry
      -- CP-element group 39: 	 branch_block_stmt_9537/assign_stmt_9563/CONCAT_u1_u16_9558_Update/$exit
      -- CP-element group 39: 	 branch_block_stmt_9537/assign_stmt_9563/CONCAT_u1_u16_9558_Update/cr
      -- CP-element group 39: 	 branch_block_stmt_9537/assign_stmt_9563/CONCAT_u1_u16_9558_Update/ca
      -- CP-element group 39: 	 branch_block_stmt_9537/assign_stmt_9563/CONCAT_u64_u128_9561_sample_start_
      -- CP-element group 39: 	 branch_block_stmt_9537/assign_stmt_9563/CONCAT_u64_u128_9561_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_9537/assign_stmt_9563/CONCAT_u64_u128_9561_update_start_
      -- CP-element group 39: 	 branch_block_stmt_9537/assign_stmt_9563/CONCAT_u64_u128_9561_update_completed_
      -- CP-element group 39: 	 branch_block_stmt_9537/assign_stmt_9563/R_Key_A_9559_sample_start_
      -- CP-element group 39: 	 branch_block_stmt_9537/assign_stmt_9563/R_Key_A_9559_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_9537/assign_stmt_9563/R_Key_A_9559_update_start_
      -- CP-element group 39: 	 branch_block_stmt_9537/assign_stmt_9563/R_Key_A_9559_update_completed_
      -- CP-element group 39: 	 branch_block_stmt_9537/assign_stmt_9563/R_Key_B_9560_sample_start_
      -- CP-element group 39: 	 branch_block_stmt_9537/assign_stmt_9563/R_Key_B_9560_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_9537/assign_stmt_9563/R_Key_B_9560_update_start_
      -- CP-element group 39: 	 branch_block_stmt_9537/assign_stmt_9563/R_Key_B_9560_update_completed_
      -- CP-element group 39: 	 branch_block_stmt_9537/assign_stmt_9563/CONCAT_u64_u128_9561_Sample/$entry
      -- CP-element group 39: 	 branch_block_stmt_9537/assign_stmt_9563/CONCAT_u64_u128_9561_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_9537/assign_stmt_9563/CONCAT_u64_u128_9561_Sample/rr
      -- CP-element group 39: 	 branch_block_stmt_9537/assign_stmt_9563/CONCAT_u64_u128_9561_Sample/ra
      -- CP-element group 39: 	 branch_block_stmt_9537/assign_stmt_9563/CONCAT_u64_u128_9561_Update/$entry
      -- CP-element group 39: 	 branch_block_stmt_9537/assign_stmt_9563/CONCAT_u64_u128_9561_Update/$exit
      -- CP-element group 39: 	 branch_block_stmt_9537/assign_stmt_9563/CONCAT_u64_u128_9561_Update/cr
      -- CP-element group 39: 	 branch_block_stmt_9537/assign_stmt_9563/CONCAT_u64_u128_9561_Update/ca
      -- CP-element group 39: 	 branch_block_stmt_9537/assign_stmt_9563/CONCAT_u16_u144_9562_Sample/$entry
      -- CP-element group 39: 	 branch_block_stmt_9537/assign_stmt_9563/CONCAT_u16_u144_9562_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_9537/assign_stmt_9563/CONCAT_u16_u144_9562_Sample/rr
      -- CP-element group 39: 	 branch_block_stmt_9537/assign_stmt_9563/CONCAT_u16_u144_9562_Sample/ra
      -- CP-element group 39: 	 branch_block_stmt_9537/assign_stmt_9563/CONCAT_u16_u144_9562_Update/$entry
      -- CP-element group 39: 	 branch_block_stmt_9537/assign_stmt_9563/CONCAT_u16_u144_9562_Update/$exit
      -- CP-element group 39: 	 branch_block_stmt_9537/assign_stmt_9563/CONCAT_u16_u144_9562_Update/cr
      -- CP-element group 39: 	 branch_block_stmt_9537/assign_stmt_9563/CONCAT_u16_u144_9562_Update/ca
      -- 
    c_block_daemon_CP_1519_elements(39) <= c_block_daemon_CP_1519_elements(22);
    -- CP-element group 40:  transition  output  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	23 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	41 
    -- CP-element group 40:  members (8) 
      -- CP-element group 40: 	 branch_block_stmt_9537/assign_stmt_9566/$entry
      -- CP-element group 40: 	 branch_block_stmt_9537/assign_stmt_9566/R_e_cmd_9565_sample_start_
      -- CP-element group 40: 	 branch_block_stmt_9537/assign_stmt_9566/R_e_cmd_9565_sample_completed_
      -- CP-element group 40: 	 branch_block_stmt_9537/assign_stmt_9566/R_e_cmd_9565_update_start_
      -- CP-element group 40: 	 branch_block_stmt_9537/assign_stmt_9566/R_e_cmd_9565_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_9537/assign_stmt_9566/WPIPE_e_cmd_pipe_9564_sample_start_
      -- CP-element group 40: 	 branch_block_stmt_9537/assign_stmt_9566/WPIPE_e_cmd_pipe_9564_Sample/$entry
      -- CP-element group 40: 	 branch_block_stmt_9537/assign_stmt_9566/WPIPE_e_cmd_pipe_9564_Sample/req
      -- 
    req_1875_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1875_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => c_block_daemon_CP_1519_elements(40), ack => WPIPE_e_cmd_pipe_9564_inst_req_0); -- 
    c_block_daemon_CP_1519_elements(40) <= c_block_daemon_CP_1519_elements(23);
    -- CP-element group 41:  transition  input  output  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	40 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	42 
    -- CP-element group 41:  members (6) 
      -- CP-element group 41: 	 branch_block_stmt_9537/assign_stmt_9566/WPIPE_e_cmd_pipe_9564_sample_completed_
      -- CP-element group 41: 	 branch_block_stmt_9537/assign_stmt_9566/WPIPE_e_cmd_pipe_9564_update_start_
      -- CP-element group 41: 	 branch_block_stmt_9537/assign_stmt_9566/WPIPE_e_cmd_pipe_9564_Sample/$exit
      -- CP-element group 41: 	 branch_block_stmt_9537/assign_stmt_9566/WPIPE_e_cmd_pipe_9564_Sample/ack
      -- CP-element group 41: 	 branch_block_stmt_9537/assign_stmt_9566/WPIPE_e_cmd_pipe_9564_Update/$entry
      -- CP-element group 41: 	 branch_block_stmt_9537/assign_stmt_9566/WPIPE_e_cmd_pipe_9564_Update/req
      -- 
    ack_1876_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_e_cmd_pipe_9564_inst_ack_0, ack => c_block_daemon_CP_1519_elements(41)); -- 
    req_1880_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1880_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => c_block_daemon_CP_1519_elements(41), ack => WPIPE_e_cmd_pipe_9564_inst_req_1); -- 
    -- CP-element group 42:  transition  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	41 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	24 
    -- CP-element group 42:  members (4) 
      -- CP-element group 42: 	 branch_block_stmt_9537/assign_stmt_9566/$exit
      -- CP-element group 42: 	 branch_block_stmt_9537/assign_stmt_9566/WPIPE_e_cmd_pipe_9564_update_completed_
      -- CP-element group 42: 	 branch_block_stmt_9537/assign_stmt_9566/WPIPE_e_cmd_pipe_9564_Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_9537/assign_stmt_9566/WPIPE_e_cmd_pipe_9564_Update/ack
      -- 
    ack_1881_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_e_cmd_pipe_9564_inst_ack_1, ack => c_block_daemon_CP_1519_elements(42)); -- 
    -- CP-element group 43:  transition  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	19 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (1) 
      -- CP-element group 43: 	 branch_block_stmt_9537/merge_stmt_9545_dead_link/$entry
      -- 
    c_block_daemon_CP_1519_elements(43) <= c_block_daemon_CP_1519_elements(19);
    -- CP-element group 44:  transition  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	19 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	46 
    -- CP-element group 44:  members (2) 
      -- CP-element group 44: 	 branch_block_stmt_9537/merge_stmt_9545__entry___PhiReq/$entry
      -- CP-element group 44: 	 branch_block_stmt_9537/merge_stmt_9545__entry___PhiReq/$exit
      -- 
    c_block_daemon_CP_1519_elements(44) <= c_block_daemon_CP_1519_elements(19);
    -- CP-element group 45:  transition  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	38 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45:  members (2) 
      -- CP-element group 45: 	 branch_block_stmt_9537/e_block_BUSY_PhiReq/$entry
      -- CP-element group 45: 	 branch_block_stmt_9537/e_block_BUSY_PhiReq/$exit
      -- 
    c_block_daemon_CP_1519_elements(45) <= c_block_daemon_CP_1519_elements(38);
    -- CP-element group 46:  merge  place  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	44 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	47 
    -- CP-element group 46:  members (1) 
      -- CP-element group 46: 	 branch_block_stmt_9537/merge_stmt_9545_PhiReqMerge
      -- 
    c_block_daemon_CP_1519_elements(46) <= OrReduce(c_block_daemon_CP_1519_elements(44) & c_block_daemon_CP_1519_elements(45));
    -- CP-element group 47:  transition  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	46 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	20 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_9537/merge_stmt_9545_PhiAck/$entry
      -- CP-element group 47: 	 branch_block_stmt_9537/merge_stmt_9545_PhiAck/$exit
      -- CP-element group 47: 	 branch_block_stmt_9537/merge_stmt_9545_PhiAck/dummy
      -- 
    c_block_daemon_CP_1519_elements(47) <= c_block_daemon_CP_1519_elements(46);
    -- CP-element group 48:  transition  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	10 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	49 
    -- CP-element group 48:  members (2) 
      -- CP-element group 48: 	 branch_block_stmt_9537/$exit
      -- CP-element group 48: 	 branch_block_stmt_9569/$entry
      -- 
    c_block_daemon_CP_1519_elements(48) <= c_block_daemon_CP_1519_elements(10);
    -- CP-element group 49:  branch  place  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	48 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	51 
    -- CP-element group 49: 	52 
    -- CP-element group 49:  members (2) 
      -- CP-element group 49: 	 branch_block_stmt_9569/branch_block_stmt_9569__entry__
      -- CP-element group 49: 	 branch_block_stmt_9569/if_stmt_9570__entry__
      -- 
    c_block_daemon_CP_1519_elements(49) <= c_block_daemon_CP_1519_elements(48);
    -- CP-element group 50:  merge  place  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	57 
    -- CP-element group 50: 	64 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	88 
    -- CP-element group 50:  members (2) 
      -- CP-element group 50: 	 branch_block_stmt_9569/branch_block_stmt_9569__exit__
      -- CP-element group 50: 	 branch_block_stmt_9569/if_stmt_9570__exit__
      -- 
    c_block_daemon_CP_1519_elements(50) <= OrReduce(c_block_daemon_CP_1519_elements(57) & c_block_daemon_CP_1519_elements(64));
    -- CP-element group 51:  transition  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	49 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (1) 
      -- CP-element group 51: 	 branch_block_stmt_9569/if_stmt_9570_dead_link/$entry
      -- 
    c_block_daemon_CP_1519_elements(51) <= c_block_daemon_CP_1519_elements(49);
    -- CP-element group 52:  transition  output  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	49 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	53 
    -- CP-element group 52:  members (17) 
      -- CP-element group 52: 	 branch_block_stmt_9569/if_stmt_9570_eval_test/branch_req
      -- CP-element group 52: 	 branch_block_stmt_9569/if_stmt_9570_eval_test/$entry
      -- CP-element group 52: 	 branch_block_stmt_9569/if_stmt_9570_eval_test/$exit
      -- CP-element group 52: 	 branch_block_stmt_9569/if_stmt_9570_eval_test/EQ_u1_u1_9573/$entry
      -- CP-element group 52: 	 branch_block_stmt_9569/if_stmt_9570_eval_test/EQ_u1_u1_9573/$exit
      -- CP-element group 52: 	 branch_block_stmt_9569/if_stmt_9570_eval_test/EQ_u1_u1_9573/EQ_u1_u1_9573_inputs/$entry
      -- CP-element group 52: 	 branch_block_stmt_9569/if_stmt_9570_eval_test/EQ_u1_u1_9573/EQ_u1_u1_9573_inputs/$exit
      -- CP-element group 52: 	 branch_block_stmt_9569/if_stmt_9570_eval_test/EQ_u1_u1_9573/SplitProtocol/$entry
      -- CP-element group 52: 	 branch_block_stmt_9569/if_stmt_9570_eval_test/EQ_u1_u1_9573/SplitProtocol/$exit
      -- CP-element group 52: 	 branch_block_stmt_9569/if_stmt_9570_eval_test/EQ_u1_u1_9573/SplitProtocol/Sample/$entry
      -- CP-element group 52: 	 branch_block_stmt_9569/if_stmt_9570_eval_test/EQ_u1_u1_9573/SplitProtocol/Sample/$exit
      -- CP-element group 52: 	 branch_block_stmt_9569/if_stmt_9570_eval_test/EQ_u1_u1_9573/SplitProtocol/Sample/rr
      -- CP-element group 52: 	 branch_block_stmt_9569/if_stmt_9570_eval_test/EQ_u1_u1_9573/SplitProtocol/Sample/ra
      -- CP-element group 52: 	 branch_block_stmt_9569/if_stmt_9570_eval_test/EQ_u1_u1_9573/SplitProtocol/Update/$entry
      -- CP-element group 52: 	 branch_block_stmt_9569/if_stmt_9570_eval_test/EQ_u1_u1_9573/SplitProtocol/Update/$exit
      -- CP-element group 52: 	 branch_block_stmt_9569/if_stmt_9570_eval_test/EQ_u1_u1_9573/SplitProtocol/Update/cr
      -- CP-element group 52: 	 branch_block_stmt_9569/if_stmt_9570_eval_test/EQ_u1_u1_9573/SplitProtocol/Update/ca
      -- 
    branch_req_1930_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1930_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => c_block_daemon_CP_1519_elements(52), ack => if_stmt_9570_branch_req_0); -- 
    c_block_daemon_CP_1519_elements(52) <= c_block_daemon_CP_1519_elements(49);
    -- CP-element group 53:  branch  place  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	52 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53: 	56 
    -- CP-element group 53:  members (1) 
      -- CP-element group 53: 	 branch_block_stmt_9569/EQ_u1_u1_9573_place
      -- 
    c_block_daemon_CP_1519_elements(53) <= c_block_daemon_CP_1519_elements(52);
    -- CP-element group 54:  transition  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	55 
    -- CP-element group 54:  members (1) 
      -- CP-element group 54: 	 branch_block_stmt_9569/if_stmt_9570_if_link/$entry
      -- 
    c_block_daemon_CP_1519_elements(54) <= c_block_daemon_CP_1519_elements(53);
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	54 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	58 
    -- CP-element group 55:  members (2) 
      -- CP-element group 55: 	 branch_block_stmt_9569/if_stmt_9570_if_link/if_choice_transition
      -- CP-element group 55: 	 branch_block_stmt_9569/if_stmt_9570_if_link/$exit
      -- 
    if_choice_transition_1935_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_9570_branch_ack_1, ack => c_block_daemon_CP_1519_elements(55)); -- 
    -- CP-element group 56:  transition  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	53 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	57 
    -- CP-element group 56:  members (1) 
      -- CP-element group 56: 	 branch_block_stmt_9569/if_stmt_9570_else_link/$entry
      -- 
    c_block_daemon_CP_1519_elements(56) <= c_block_daemon_CP_1519_elements(53);
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	56 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	50 
    -- CP-element group 57:  members (2) 
      -- CP-element group 57: 	 branch_block_stmt_9569/if_stmt_9570_else_link/else_choice_transition
      -- CP-element group 57: 	 branch_block_stmt_9569/if_stmt_9570_else_link/$exit
      -- 
    else_choice_transition_1939_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_9570_branch_ack_0, ack => c_block_daemon_CP_1519_elements(57)); -- 
    -- CP-element group 58:  place  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	55 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	65 
    -- CP-element group 58:  members (1) 
      -- CP-element group 58: 	 branch_block_stmt_9569/assign_stmt_9576__entry__
      -- 
    c_block_daemon_CP_1519_elements(58) <= c_block_daemon_CP_1519_elements(55);
    -- CP-element group 59:  branch  place  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	67 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	83 
    -- CP-element group 59: 	84 
    -- CP-element group 59:  members (2) 
      -- CP-element group 59: 	 branch_block_stmt_9569/merge_stmt_9577__entry__
      -- CP-element group 59: 	 branch_block_stmt_9569/assign_stmt_9576__exit__
      -- 
    c_block_daemon_CP_1519_elements(59) <= c_block_daemon_CP_1519_elements(67);
    -- CP-element group 60:  merge  place  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	87 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	68 
    -- CP-element group 60:  members (2) 
      -- CP-element group 60: 	 branch_block_stmt_9569/assign_stmt_9580__entry__
      -- CP-element group 60: 	 branch_block_stmt_9569/merge_stmt_9577__exit__
      -- 
    c_block_daemon_CP_1519_elements(60) <= c_block_daemon_CP_1519_elements(87);
    -- CP-element group 61:  branch  place  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	70 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	71 
    -- CP-element group 61: 	72 
    -- CP-element group 61:  members (2) 
      -- CP-element group 61: 	 branch_block_stmt_9569/if_stmt_9581__entry__
      -- CP-element group 61: 	 branch_block_stmt_9569/assign_stmt_9580__exit__
      -- 
    c_block_daemon_CP_1519_elements(61) <= c_block_daemon_CP_1519_elements(70);
    -- CP-element group 62:  merge  place  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	77 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	79 
    -- CP-element group 62:  members (2) 
      -- CP-element group 62: 	 branch_block_stmt_9569/if_stmt_9581__exit__
      -- CP-element group 62: 	 branch_block_stmt_9569/assign_stmt_9595__entry__
      -- 
    c_block_daemon_CP_1519_elements(62) <= c_block_daemon_CP_1519_elements(77);
    -- CP-element group 63:  place  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	79 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	80 
    -- CP-element group 63:  members (2) 
      -- CP-element group 63: 	 branch_block_stmt_9569/assign_stmt_9595__exit__
      -- CP-element group 63: 	 branch_block_stmt_9569/assign_stmt_9598__entry__
      -- 
    c_block_daemon_CP_1519_elements(63) <= c_block_daemon_CP_1519_elements(79);
    -- CP-element group 64:  place  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	82 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	50 
    -- CP-element group 64:  members (1) 
      -- CP-element group 64: 	 branch_block_stmt_9569/assign_stmt_9598__exit__
      -- 
    c_block_daemon_CP_1519_elements(64) <= c_block_daemon_CP_1519_elements(82);
    -- CP-element group 65:  transition  output  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	58 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	66 
    -- CP-element group 65:  members (4) 
      -- CP-element group 65: 	 branch_block_stmt_9569/assign_stmt_9576/WPIPE_status_out_9574_sample_start_
      -- CP-element group 65: 	 branch_block_stmt_9569/assign_stmt_9576/WPIPE_status_out_9574_Sample/req
      -- CP-element group 65: 	 branch_block_stmt_9569/assign_stmt_9576/$entry
      -- CP-element group 65: 	 branch_block_stmt_9569/assign_stmt_9576/WPIPE_status_out_9574_Sample/$entry
      -- 
    req_1962_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1962_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => c_block_daemon_CP_1519_elements(65), ack => WPIPE_status_out_9574_inst_req_0); -- 
    c_block_daemon_CP_1519_elements(65) <= c_block_daemon_CP_1519_elements(58);
    -- CP-element group 66:  transition  input  output  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	65 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66:  members (6) 
      -- CP-element group 66: 	 branch_block_stmt_9569/assign_stmt_9576/WPIPE_status_out_9574_update_start_
      -- CP-element group 66: 	 branch_block_stmt_9569/assign_stmt_9576/WPIPE_status_out_9574_sample_completed_
      -- CP-element group 66: 	 branch_block_stmt_9569/assign_stmt_9576/WPIPE_status_out_9574_Update/req
      -- CP-element group 66: 	 branch_block_stmt_9569/assign_stmt_9576/WPIPE_status_out_9574_Update/$entry
      -- CP-element group 66: 	 branch_block_stmt_9569/assign_stmt_9576/WPIPE_status_out_9574_Sample/ack
      -- CP-element group 66: 	 branch_block_stmt_9569/assign_stmt_9576/WPIPE_status_out_9574_Sample/$exit
      -- 
    ack_1963_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_status_out_9574_inst_ack_0, ack => c_block_daemon_CP_1519_elements(66)); -- 
    req_1967_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1967_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => c_block_daemon_CP_1519_elements(66), ack => WPIPE_status_out_9574_inst_req_1); -- 
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	59 
    -- CP-element group 67:  members (4) 
      -- CP-element group 67: 	 branch_block_stmt_9569/assign_stmt_9576/$exit
      -- CP-element group 67: 	 branch_block_stmt_9569/assign_stmt_9576/WPIPE_status_out_9574_Update/ack
      -- CP-element group 67: 	 branch_block_stmt_9569/assign_stmt_9576/WPIPE_status_out_9574_Update/$exit
      -- CP-element group 67: 	 branch_block_stmt_9569/assign_stmt_9576/WPIPE_status_out_9574_update_completed_
      -- 
    ack_1968_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_status_out_9574_inst_ack_1, ack => c_block_daemon_CP_1519_elements(67)); -- 
    -- CP-element group 68:  transition  output  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	60 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	69 
    -- CP-element group 68:  members (4) 
      -- CP-element group 68: 	 branch_block_stmt_9569/assign_stmt_9580/RPIPE_d_block_done_9579_Sample/$entry
      -- CP-element group 68: 	 branch_block_stmt_9569/assign_stmt_9580/RPIPE_d_block_done_9579_sample_start_
      -- CP-element group 68: 	 branch_block_stmt_9569/assign_stmt_9580/RPIPE_d_block_done_9579_Sample/rr
      -- CP-element group 68: 	 branch_block_stmt_9569/assign_stmt_9580/$entry
      -- 
    rr_1979_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1979_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => c_block_daemon_CP_1519_elements(68), ack => RPIPE_d_block_done_9579_inst_req_0); -- 
    c_block_daemon_CP_1519_elements(68) <= c_block_daemon_CP_1519_elements(60);
    -- CP-element group 69:  transition  input  output  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	68 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	70 
    -- CP-element group 69:  members (6) 
      -- CP-element group 69: 	 branch_block_stmt_9569/assign_stmt_9580/RPIPE_d_block_done_9579_Update/cr
      -- CP-element group 69: 	 branch_block_stmt_9569/assign_stmt_9580/RPIPE_d_block_done_9579_Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_9569/assign_stmt_9580/RPIPE_d_block_done_9579_Sample/ra
      -- CP-element group 69: 	 branch_block_stmt_9569/assign_stmt_9580/RPIPE_d_block_done_9579_update_start_
      -- CP-element group 69: 	 branch_block_stmt_9569/assign_stmt_9580/RPIPE_d_block_done_9579_sample_completed_
      -- CP-element group 69: 	 branch_block_stmt_9569/assign_stmt_9580/RPIPE_d_block_done_9579_Sample/$exit
      -- 
    ra_1980_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_d_block_done_9579_inst_ack_0, ack => c_block_daemon_CP_1519_elements(69)); -- 
    cr_1984_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1984_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => c_block_daemon_CP_1519_elements(69), ack => RPIPE_d_block_done_9579_inst_req_1); -- 
    -- CP-element group 70:  transition  input  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	69 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	61 
    -- CP-element group 70:  members (4) 
      -- CP-element group 70: 	 branch_block_stmt_9569/assign_stmt_9580/RPIPE_d_block_done_9579_Update/$exit
      -- CP-element group 70: 	 branch_block_stmt_9569/assign_stmt_9580/RPIPE_d_block_done_9579_Update/ca
      -- CP-element group 70: 	 branch_block_stmt_9569/assign_stmt_9580/RPIPE_d_block_done_9579_update_completed_
      -- CP-element group 70: 	 branch_block_stmt_9569/assign_stmt_9580/$exit
      -- 
    ca_1985_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_d_block_done_9579_inst_ack_1, ack => c_block_daemon_CP_1519_elements(70)); -- 
    -- CP-element group 71:  transition  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	61 
    -- CP-element group 71: successors 
    -- CP-element group 71:  members (1) 
      -- CP-element group 71: 	 branch_block_stmt_9569/if_stmt_9581_dead_link/$entry
      -- 
    c_block_daemon_CP_1519_elements(71) <= c_block_daemon_CP_1519_elements(61);
    -- CP-element group 72:  transition  output  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	61 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	73 
    -- CP-element group 72:  members (17) 
      -- CP-element group 72: 	 branch_block_stmt_9569/if_stmt_9581_eval_test/EQ_u1_u1_9584/SplitProtocol/$entry
      -- CP-element group 72: 	 branch_block_stmt_9569/if_stmt_9581_eval_test/EQ_u1_u1_9584/SplitProtocol/$exit
      -- CP-element group 72: 	 branch_block_stmt_9569/if_stmt_9581_eval_test/EQ_u1_u1_9584/EQ_u1_u1_9584_inputs/$entry
      -- CP-element group 72: 	 branch_block_stmt_9569/if_stmt_9581_eval_test/EQ_u1_u1_9584/EQ_u1_u1_9584_inputs/$exit
      -- CP-element group 72: 	 branch_block_stmt_9569/if_stmt_9581_eval_test/branch_req
      -- CP-element group 72: 	 branch_block_stmt_9569/if_stmt_9581_eval_test/EQ_u1_u1_9584/SplitProtocol/Sample/rr
      -- CP-element group 72: 	 branch_block_stmt_9569/if_stmt_9581_eval_test/EQ_u1_u1_9584/SplitProtocol/Sample/ra
      -- CP-element group 72: 	 branch_block_stmt_9569/if_stmt_9581_eval_test/EQ_u1_u1_9584/SplitProtocol/Update/cr
      -- CP-element group 72: 	 branch_block_stmt_9569/if_stmt_9581_eval_test/EQ_u1_u1_9584/SplitProtocol/Update/ca
      -- CP-element group 72: 	 branch_block_stmt_9569/if_stmt_9581_eval_test/$entry
      -- CP-element group 72: 	 branch_block_stmt_9569/if_stmt_9581_eval_test/$exit
      -- CP-element group 72: 	 branch_block_stmt_9569/if_stmt_9581_eval_test/EQ_u1_u1_9584/$entry
      -- CP-element group 72: 	 branch_block_stmt_9569/if_stmt_9581_eval_test/EQ_u1_u1_9584/$exit
      -- CP-element group 72: 	 branch_block_stmt_9569/if_stmt_9581_eval_test/EQ_u1_u1_9584/SplitProtocol/Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_9569/if_stmt_9581_eval_test/EQ_u1_u1_9584/SplitProtocol/Sample/$exit
      -- CP-element group 72: 	 branch_block_stmt_9569/if_stmt_9581_eval_test/EQ_u1_u1_9584/SplitProtocol/Update/$entry
      -- CP-element group 72: 	 branch_block_stmt_9569/if_stmt_9581_eval_test/EQ_u1_u1_9584/SplitProtocol/Update/$exit
      -- 
    branch_req_2012_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2012_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => c_block_daemon_CP_1519_elements(72), ack => if_stmt_9581_branch_req_0); -- 
    c_block_daemon_CP_1519_elements(72) <= c_block_daemon_CP_1519_elements(61);
    -- CP-element group 73:  branch  place  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	72 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	74 
    -- CP-element group 73: 	76 
    -- CP-element group 73:  members (1) 
      -- CP-element group 73: 	 branch_block_stmt_9569/EQ_u1_u1_9584_place
      -- 
    c_block_daemon_CP_1519_elements(73) <= c_block_daemon_CP_1519_elements(72);
    -- CP-element group 74:  transition  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	73 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	75 
    -- CP-element group 74:  members (1) 
      -- CP-element group 74: 	 branch_block_stmt_9569/if_stmt_9581_if_link/$entry
      -- 
    c_block_daemon_CP_1519_elements(74) <= c_block_daemon_CP_1519_elements(73);
    -- CP-element group 75:  transition  input  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	74 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	78 
    -- CP-element group 75:  members (2) 
      -- CP-element group 75: 	 branch_block_stmt_9569/if_stmt_9581_if_link/$exit
      -- CP-element group 75: 	 branch_block_stmt_9569/if_stmt_9581_if_link/if_choice_transition
      -- 
    if_choice_transition_2017_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_9581_branch_ack_1, ack => c_block_daemon_CP_1519_elements(75)); -- 
    -- CP-element group 76:  transition  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	73 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	77 
    -- CP-element group 76:  members (1) 
      -- CP-element group 76: 	 branch_block_stmt_9569/if_stmt_9581_else_link/$entry
      -- 
    c_block_daemon_CP_1519_elements(76) <= c_block_daemon_CP_1519_elements(73);
    -- CP-element group 77:  transition  input  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	76 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	62 
    -- CP-element group 77:  members (2) 
      -- CP-element group 77: 	 branch_block_stmt_9569/if_stmt_9581_else_link/$exit
      -- CP-element group 77: 	 branch_block_stmt_9569/if_stmt_9581_else_link/else_choice_transition
      -- 
    else_choice_transition_2021_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_9581_branch_ack_0, ack => c_block_daemon_CP_1519_elements(77)); -- 
    -- CP-element group 78:  place  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	75 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	85 
    -- CP-element group 78:  members (1) 
      -- CP-element group 78: 	 branch_block_stmt_9569/d_block_BUSY
      -- 
    c_block_daemon_CP_1519_elements(78) <= c_block_daemon_CP_1519_elements(75);
    -- CP-element group 79:  join  fork  transition  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	62 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	63 
    -- CP-element group 79:  members (54) 
      -- CP-element group 79: 	 branch_block_stmt_9569/assign_stmt_9595/R_got_new_key_9588_sample_completed_
      -- CP-element group 79: 	 branch_block_stmt_9569/assign_stmt_9595/R_got_new_key_9588_update_start_
      -- CP-element group 79: 	 branch_block_stmt_9569/assign_stmt_9595/R_got_new_key_9588_update_completed_
      -- CP-element group 79: 	 branch_block_stmt_9569/assign_stmt_9595/$exit
      -- CP-element group 79: 	 branch_block_stmt_9569/assign_stmt_9595/R_Key_B_9592_update_completed_
      -- CP-element group 79: 	 branch_block_stmt_9569/assign_stmt_9595/CONCAT_u64_u128_9593_Sample/$entry
      -- CP-element group 79: 	 branch_block_stmt_9569/assign_stmt_9595/CONCAT_u64_u128_9593_Sample/$exit
      -- CP-element group 79: 	 branch_block_stmt_9569/assign_stmt_9595/CONCAT_u64_u128_9593_Sample/rr
      -- CP-element group 79: 	 branch_block_stmt_9569/assign_stmt_9595/CONCAT_u64_u128_9593_Sample/ra
      -- CP-element group 79: 	 branch_block_stmt_9569/assign_stmt_9595/CONCAT_u1_u16_9590_Update/cr
      -- CP-element group 79: 	 branch_block_stmt_9569/assign_stmt_9595/CONCAT_u1_u16_9590_Update/ca
      -- CP-element group 79: 	 branch_block_stmt_9569/assign_stmt_9595/CONCAT_u64_u128_9593_sample_start_
      -- CP-element group 79: 	 branch_block_stmt_9569/assign_stmt_9595/CONCAT_u64_u128_9593_sample_completed_
      -- CP-element group 79: 	 branch_block_stmt_9569/assign_stmt_9595/CONCAT_u64_u128_9593_update_start_
      -- CP-element group 79: 	 branch_block_stmt_9569/assign_stmt_9595/CONCAT_u64_u128_9593_update_completed_
      -- CP-element group 79: 	 branch_block_stmt_9569/assign_stmt_9595/R_Key_A_9591_sample_start_
      -- CP-element group 79: 	 branch_block_stmt_9569/assign_stmt_9595/CONCAT_u1_u16_9590_Sample/$entry
      -- CP-element group 79: 	 branch_block_stmt_9569/assign_stmt_9595/CONCAT_u1_u16_9590_Sample/$exit
      -- CP-element group 79: 	 branch_block_stmt_9569/assign_stmt_9595/CONCAT_u1_u16_9590_Sample/rr
      -- CP-element group 79: 	 branch_block_stmt_9569/assign_stmt_9595/CONCAT_u1_u16_9590_Sample/ra
      -- CP-element group 79: 	 branch_block_stmt_9569/assign_stmt_9595/CONCAT_u1_u16_9590_Update/$entry
      -- CP-element group 79: 	 branch_block_stmt_9569/assign_stmt_9595/CONCAT_u1_u16_9590_Update/$exit
      -- CP-element group 79: 	 branch_block_stmt_9569/assign_stmt_9595/R_Key_A_9591_sample_completed_
      -- CP-element group 79: 	 branch_block_stmt_9569/assign_stmt_9595/R_Key_A_9591_update_start_
      -- CP-element group 79: 	 branch_block_stmt_9569/assign_stmt_9595/R_Key_A_9591_update_completed_
      -- CP-element group 79: 	 branch_block_stmt_9569/assign_stmt_9595/R_Key_B_9592_sample_start_
      -- CP-element group 79: 	 branch_block_stmt_9569/assign_stmt_9595/R_Key_B_9592_sample_completed_
      -- CP-element group 79: 	 branch_block_stmt_9569/assign_stmt_9595/R_Key_B_9592_update_start_
      -- CP-element group 79: 	 branch_block_stmt_9569/assign_stmt_9595/CONCAT_u1_u16_9590_update_start_
      -- CP-element group 79: 	 branch_block_stmt_9569/assign_stmt_9595/CONCAT_u1_u16_9590_update_completed_
      -- CP-element group 79: 	 branch_block_stmt_9569/assign_stmt_9595/R_got_new_key_9588_sample_start_
      -- CP-element group 79: 	 branch_block_stmt_9569/assign_stmt_9595/R_count_9589_sample_start_
      -- CP-element group 79: 	 branch_block_stmt_9569/assign_stmt_9595/R_count_9589_sample_completed_
      -- CP-element group 79: 	 branch_block_stmt_9569/assign_stmt_9595/R_count_9589_update_start_
      -- CP-element group 79: 	 branch_block_stmt_9569/assign_stmt_9595/R_count_9589_update_completed_
      -- CP-element group 79: 	 branch_block_stmt_9569/assign_stmt_9595/CONCAT_u16_u144_9594_sample_start_
      -- CP-element group 79: 	 branch_block_stmt_9569/assign_stmt_9595/CONCAT_u16_u144_9594_sample_completed_
      -- CP-element group 79: 	 branch_block_stmt_9569/assign_stmt_9595/CONCAT_u16_u144_9594_update_start_
      -- CP-element group 79: 	 branch_block_stmt_9569/assign_stmt_9595/$entry
      -- CP-element group 79: 	 branch_block_stmt_9569/assign_stmt_9595/CONCAT_u16_u144_9594_update_completed_
      -- CP-element group 79: 	 branch_block_stmt_9569/assign_stmt_9595/CONCAT_u1_u16_9590_sample_start_
      -- CP-element group 79: 	 branch_block_stmt_9569/assign_stmt_9595/CONCAT_u1_u16_9590_sample_completed_
      -- CP-element group 79: 	 branch_block_stmt_9569/assign_stmt_9595/CONCAT_u64_u128_9593_Update/$entry
      -- CP-element group 79: 	 branch_block_stmt_9569/assign_stmt_9595/CONCAT_u64_u128_9593_Update/$exit
      -- CP-element group 79: 	 branch_block_stmt_9569/assign_stmt_9595/CONCAT_u64_u128_9593_Update/cr
      -- CP-element group 79: 	 branch_block_stmt_9569/assign_stmt_9595/CONCAT_u64_u128_9593_Update/ca
      -- CP-element group 79: 	 branch_block_stmt_9569/assign_stmt_9595/CONCAT_u16_u144_9594_Sample/$entry
      -- CP-element group 79: 	 branch_block_stmt_9569/assign_stmt_9595/CONCAT_u16_u144_9594_Sample/$exit
      -- CP-element group 79: 	 branch_block_stmt_9569/assign_stmt_9595/CONCAT_u16_u144_9594_Sample/rr
      -- CP-element group 79: 	 branch_block_stmt_9569/assign_stmt_9595/CONCAT_u16_u144_9594_Sample/ra
      -- CP-element group 79: 	 branch_block_stmt_9569/assign_stmt_9595/CONCAT_u16_u144_9594_Update/$entry
      -- CP-element group 79: 	 branch_block_stmt_9569/assign_stmt_9595/CONCAT_u16_u144_9594_Update/$exit
      -- CP-element group 79: 	 branch_block_stmt_9569/assign_stmt_9595/CONCAT_u16_u144_9594_Update/cr
      -- CP-element group 79: 	 branch_block_stmt_9569/assign_stmt_9595/CONCAT_u16_u144_9594_Update/ca
      -- 
    c_block_daemon_CP_1519_elements(79) <= c_block_daemon_CP_1519_elements(62);
    -- CP-element group 80:  transition  output  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	63 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	81 
    -- CP-element group 80:  members (8) 
      -- CP-element group 80: 	 branch_block_stmt_9569/assign_stmt_9598/$entry
      -- CP-element group 80: 	 branch_block_stmt_9569/assign_stmt_9598/R_d_cmd_9597_sample_start_
      -- CP-element group 80: 	 branch_block_stmt_9569/assign_stmt_9598/R_d_cmd_9597_sample_completed_
      -- CP-element group 80: 	 branch_block_stmt_9569/assign_stmt_9598/R_d_cmd_9597_update_start_
      -- CP-element group 80: 	 branch_block_stmt_9569/assign_stmt_9598/R_d_cmd_9597_update_completed_
      -- CP-element group 80: 	 branch_block_stmt_9569/assign_stmt_9598/WPIPE_d_cmd_pipe_9596_sample_start_
      -- CP-element group 80: 	 branch_block_stmt_9569/assign_stmt_9598/WPIPE_d_cmd_pipe_9596_Sample/$entry
      -- CP-element group 80: 	 branch_block_stmt_9569/assign_stmt_9598/WPIPE_d_cmd_pipe_9596_Sample/req
      -- 
    req_2098_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2098_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => c_block_daemon_CP_1519_elements(80), ack => WPIPE_d_cmd_pipe_9596_inst_req_0); -- 
    c_block_daemon_CP_1519_elements(80) <= c_block_daemon_CP_1519_elements(63);
    -- CP-element group 81:  transition  input  output  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	80 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	82 
    -- CP-element group 81:  members (6) 
      -- CP-element group 81: 	 branch_block_stmt_9569/assign_stmt_9598/WPIPE_d_cmd_pipe_9596_sample_completed_
      -- CP-element group 81: 	 branch_block_stmt_9569/assign_stmt_9598/WPIPE_d_cmd_pipe_9596_update_start_
      -- CP-element group 81: 	 branch_block_stmt_9569/assign_stmt_9598/WPIPE_d_cmd_pipe_9596_Sample/$exit
      -- CP-element group 81: 	 branch_block_stmt_9569/assign_stmt_9598/WPIPE_d_cmd_pipe_9596_Sample/ack
      -- CP-element group 81: 	 branch_block_stmt_9569/assign_stmt_9598/WPIPE_d_cmd_pipe_9596_Update/$entry
      -- CP-element group 81: 	 branch_block_stmt_9569/assign_stmt_9598/WPIPE_d_cmd_pipe_9596_Update/req
      -- 
    ack_2099_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_d_cmd_pipe_9596_inst_ack_0, ack => c_block_daemon_CP_1519_elements(81)); -- 
    req_2103_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2103_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => c_block_daemon_CP_1519_elements(81), ack => WPIPE_d_cmd_pipe_9596_inst_req_1); -- 
    -- CP-element group 82:  transition  input  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	81 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	64 
    -- CP-element group 82:  members (4) 
      -- CP-element group 82: 	 branch_block_stmt_9569/assign_stmt_9598/$exit
      -- CP-element group 82: 	 branch_block_stmt_9569/assign_stmt_9598/WPIPE_d_cmd_pipe_9596_update_completed_
      -- CP-element group 82: 	 branch_block_stmt_9569/assign_stmt_9598/WPIPE_d_cmd_pipe_9596_Update/$exit
      -- CP-element group 82: 	 branch_block_stmt_9569/assign_stmt_9598/WPIPE_d_cmd_pipe_9596_Update/ack
      -- 
    ack_2104_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_d_cmd_pipe_9596_inst_ack_1, ack => c_block_daemon_CP_1519_elements(82)); -- 
    -- CP-element group 83:  transition  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	59 
    -- CP-element group 83: successors 
    -- CP-element group 83:  members (1) 
      -- CP-element group 83: 	 branch_block_stmt_9569/merge_stmt_9577_dead_link/$entry
      -- 
    c_block_daemon_CP_1519_elements(83) <= c_block_daemon_CP_1519_elements(59);
    -- CP-element group 84:  transition  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	59 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	86 
    -- CP-element group 84:  members (2) 
      -- CP-element group 84: 	 branch_block_stmt_9569/merge_stmt_9577__entry___PhiReq/$entry
      -- CP-element group 84: 	 branch_block_stmt_9569/merge_stmt_9577__entry___PhiReq/$exit
      -- 
    c_block_daemon_CP_1519_elements(84) <= c_block_daemon_CP_1519_elements(59);
    -- CP-element group 85:  transition  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	78 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	86 
    -- CP-element group 85:  members (2) 
      -- CP-element group 85: 	 branch_block_stmt_9569/d_block_BUSY_PhiReq/$entry
      -- CP-element group 85: 	 branch_block_stmt_9569/d_block_BUSY_PhiReq/$exit
      -- 
    c_block_daemon_CP_1519_elements(85) <= c_block_daemon_CP_1519_elements(78);
    -- CP-element group 86:  merge  place  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	84 
    -- CP-element group 86: 	85 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	87 
    -- CP-element group 86:  members (1) 
      -- CP-element group 86: 	 branch_block_stmt_9569/merge_stmt_9577_PhiReqMerge
      -- 
    c_block_daemon_CP_1519_elements(86) <= OrReduce(c_block_daemon_CP_1519_elements(84) & c_block_daemon_CP_1519_elements(85));
    -- CP-element group 87:  transition  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	86 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	60 
    -- CP-element group 87:  members (3) 
      -- CP-element group 87: 	 branch_block_stmt_9569/merge_stmt_9577_PhiAck/$entry
      -- CP-element group 87: 	 branch_block_stmt_9569/merge_stmt_9577_PhiAck/$exit
      -- CP-element group 87: 	 branch_block_stmt_9569/merge_stmt_9577_PhiAck/dummy
      -- 
    c_block_daemon_CP_1519_elements(87) <= c_block_daemon_CP_1519_elements(86);
    -- CP-element group 88:  transition  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	50 
    -- CP-element group 88: successors 
    -- CP-element group 88:  members (2) 
      -- CP-element group 88: 	 $exit
      -- CP-element group 88: 	 branch_block_stmt_9569/$exit
      -- 
    c_block_daemon_CP_1519_elements(88) <= c_block_daemon_CP_1519_elements(50);
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal CONCAT_u1_u16_9558_wire : std_logic_vector(15 downto 0);
    signal CONCAT_u1_u16_9590_wire : std_logic_vector(15 downto 0);
    signal CONCAT_u64_u128_9561_wire : std_logic_vector(127 downto 0);
    signal CONCAT_u64_u128_9593_wire : std_logic_vector(127 downto 0);
    signal ED_9512 : std_logic_vector(0 downto 0);
    signal EQ_u1_u1_9541_wire : std_logic_vector(0 downto 0);
    signal EQ_u1_u1_9552_wire : std_logic_vector(0 downto 0);
    signal EQ_u1_u1_9573_wire : std_logic_vector(0 downto 0);
    signal EQ_u1_u1_9584_wire : std_logic_vector(0 downto 0);
    signal Key_A_9531 : std_logic_vector(63 downto 0);
    signal Key_B_9535 : std_logic_vector(63 downto 0);
    signal command_9508 : std_logic_vector(63 downto 0);
    signal count_9528 : std_logic_vector(14 downto 0);
    signal d_cmd_9595 : std_logic_vector(143 downto 0);
    signal d_status_9580 : std_logic_vector(0 downto 0);
    signal e_cmd_9563 : std_logic_vector(143 downto 0);
    signal e_status_9548 : std_logic_vector(0 downto 0);
    signal got_new_key_9520 : std_logic_vector(0 downto 0);
    signal konst_9540_wire_constant : std_logic_vector(0 downto 0);
    signal konst_9543_wire_constant : std_logic_vector(63 downto 0);
    signal konst_9551_wire_constant : std_logic_vector(0 downto 0);
    signal konst_9572_wire_constant : std_logic_vector(0 downto 0);
    signal konst_9575_wire_constant : std_logic_vector(63 downto 0);
    signal konst_9583_wire_constant : std_logic_vector(0 downto 0);
    signal mode_9516 : std_logic_vector(2 downto 0);
    signal unused_44_9524 : std_logic_vector(43 downto 0);
    -- 
  begin -- 
    konst_9540_wire_constant <= "0";
    konst_9543_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    konst_9551_wire_constant <= "0";
    konst_9572_wire_constant <= "1";
    konst_9575_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    konst_9583_wire_constant <= "0";
    -- flow-through slice operator slice_9511_inst
    ED_9512 <= command_9508(63 downto 63);
    -- flow-through slice operator slice_9515_inst
    mode_9516 <= command_9508(62 downto 60);
    -- flow-through slice operator slice_9519_inst
    got_new_key_9520 <= command_9508(59 downto 59);
    -- flow-through slice operator slice_9523_inst
    unused_44_9524 <= command_9508(58 downto 15);
    -- flow-through slice operator slice_9527_inst
    count_9528 <= command_9508(14 downto 0);
    if_stmt_9538_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= EQ_u1_u1_9541_wire;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_9538_branch", condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_9538_branch_req_0,
          ack0 => if_stmt_9538_branch_ack_0,
          ack1 => if_stmt_9538_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_9549_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= EQ_u1_u1_9552_wire;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_9549_branch", condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_9549_branch_req_0,
          ack0 => if_stmt_9549_branch_ack_0,
          ack1 => if_stmt_9549_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_9570_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= EQ_u1_u1_9573_wire;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_9570_branch", condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_9570_branch_req_0,
          ack0 => if_stmt_9570_branch_ack_0,
          ack1 => if_stmt_9570_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_9581_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= EQ_u1_u1_9584_wire;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_9581_branch", condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_9581_branch_req_0,
          ack0 => if_stmt_9581_branch_ack_0,
          ack1 => if_stmt_9581_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator CONCAT_u16_u144_9562_inst
    process(CONCAT_u1_u16_9558_wire, CONCAT_u64_u128_9561_wire) -- 
      variable tmp_var : std_logic_vector(143 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u1_u16_9558_wire, CONCAT_u64_u128_9561_wire, tmp_var);
      e_cmd_9563 <= tmp_var; -- 
    end process;
    -- binary operator CONCAT_u16_u144_9594_inst
    process(CONCAT_u1_u16_9590_wire, CONCAT_u64_u128_9593_wire) -- 
      variable tmp_var : std_logic_vector(143 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u1_u16_9590_wire, CONCAT_u64_u128_9593_wire, tmp_var);
      d_cmd_9595 <= tmp_var; -- 
    end process;
    -- binary operator CONCAT_u1_u16_9558_inst
    process(got_new_key_9520, count_9528) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApConcat_proc(got_new_key_9520, count_9528, tmp_var);
      CONCAT_u1_u16_9558_wire <= tmp_var; -- 
    end process;
    -- binary operator CONCAT_u1_u16_9590_inst
    process(got_new_key_9520, count_9528) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApConcat_proc(got_new_key_9520, count_9528, tmp_var);
      CONCAT_u1_u16_9590_wire <= tmp_var; -- 
    end process;
    -- binary operator CONCAT_u64_u128_9561_inst
    process(Key_A_9531, Key_B_9535) -- 
      variable tmp_var : std_logic_vector(127 downto 0); -- 
    begin -- 
      ApConcat_proc(Key_A_9531, Key_B_9535, tmp_var);
      CONCAT_u64_u128_9561_wire <= tmp_var; -- 
    end process;
    -- binary operator CONCAT_u64_u128_9593_inst
    process(Key_A_9531, Key_B_9535) -- 
      variable tmp_var : std_logic_vector(127 downto 0); -- 
    begin -- 
      ApConcat_proc(Key_A_9531, Key_B_9535, tmp_var);
      CONCAT_u64_u128_9593_wire <= tmp_var; -- 
    end process;
    -- binary operator EQ_u1_u1_9541_inst
    process(ED_9512) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(ED_9512, konst_9540_wire_constant, tmp_var);
      EQ_u1_u1_9541_wire <= tmp_var; -- 
    end process;
    -- binary operator EQ_u1_u1_9552_inst
    process(e_status_9548) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(e_status_9548, konst_9551_wire_constant, tmp_var);
      EQ_u1_u1_9552_wire <= tmp_var; -- 
    end process;
    -- binary operator EQ_u1_u1_9573_inst
    process(ED_9512) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(ED_9512, konst_9572_wire_constant, tmp_var);
      EQ_u1_u1_9573_wire <= tmp_var; -- 
    end process;
    -- binary operator EQ_u1_u1_9584_inst
    process(d_status_9580) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(d_status_9580, konst_9583_wire_constant, tmp_var);
      EQ_u1_u1_9584_wire <= tmp_var; -- 
    end process;
    -- shared inport operator group (0) : RPIPE_cmd_in_9507_inst RPIPE_cmd_in_9530_inst RPIPE_cmd_in_9534_inst 
    InportGroup0: Block -- 
      signal data_out: std_logic_vector(191 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 2 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 2 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 2 downto 0);
      signal guard_vector : std_logic_vector( 2 downto 0);
      constant outBUFs : IntegerArray(2 downto 0) := (2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(2 downto 0) := (0 => true, 1 => true, 2 => false);
      constant guardBuffering: IntegerArray(2 downto 0)  := (0 => 2, 1 => 2, 2 => 2);
      -- 
    begin -- 
      reqL_unguarded(2) <= RPIPE_cmd_in_9507_inst_req_0;
      reqL_unguarded(1) <= RPIPE_cmd_in_9530_inst_req_0;
      reqL_unguarded(0) <= RPIPE_cmd_in_9534_inst_req_0;
      RPIPE_cmd_in_9507_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_cmd_in_9530_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_cmd_in_9534_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(2) <= RPIPE_cmd_in_9507_inst_req_1;
      reqR_unguarded(1) <= RPIPE_cmd_in_9530_inst_req_1;
      reqR_unguarded(0) <= RPIPE_cmd_in_9534_inst_req_1;
      RPIPE_cmd_in_9507_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_cmd_in_9530_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_cmd_in_9534_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= got_new_key_9520(0);
      guard_vector(1)  <= got_new_key_9520(0);
      guard_vector(2)  <=  '1';
      gI: SplitGuardInterface generic map(name => "gI", nreqs => 3, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      command_9508 <= data_out(191 downto 128);
      Key_A_9531 <= data_out(127 downto 64);
      Key_B_9535 <= data_out(63 downto 0);
      cmd_in_read_0: InputPortRevised -- 
        generic map ( name => "cmd_in_read_0", data_width => 64,  num_reqs => 3,  output_buffering => outBUFs,   no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => cmd_in_pipe_read_req(0),
          oack => cmd_in_pipe_read_ack(0),
          odata => cmd_in_pipe_read_data(63 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared inport operator group (1) : RPIPE_d_block_done_9579_inst 
    InportGroup1: Block -- 
      signal data_out: std_logic_vector(0 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_d_block_done_9579_inst_req_0;
      RPIPE_d_block_done_9579_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_d_block_done_9579_inst_req_1;
      RPIPE_d_block_done_9579_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      gI: SplitGuardInterface generic map(name => "gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      d_status_9580 <= data_out(0 downto 0);
      d_block_done_read_1: InputPortRevised -- 
        generic map ( name => "d_block_done_read_1", data_width => 1,  num_reqs => 1,  output_buffering => outBUFs,   no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => d_block_done_pipe_read_req(0),
          oack => d_block_done_pipe_read_ack(0),
          odata => d_block_done_pipe_read_data(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 1
    -- shared inport operator group (2) : RPIPE_e_block_done_9547_inst 
    InportGroup2: Block -- 
      signal data_out: std_logic_vector(0 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_e_block_done_9547_inst_req_0;
      RPIPE_e_block_done_9547_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_e_block_done_9547_inst_req_1;
      RPIPE_e_block_done_9547_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      gI: SplitGuardInterface generic map(name => "gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      e_status_9548 <= data_out(0 downto 0);
      e_block_done_read_2: InputPortRevised -- 
        generic map ( name => "e_block_done_read_2", data_width => 1,  num_reqs => 1,  output_buffering => outBUFs,   no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => e_block_done_pipe_read_req(0),
          oack => e_block_done_pipe_read_ack(0),
          odata => e_block_done_pipe_read_data(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 2
    -- shared outport operator group (0) : WPIPE_d_cmd_pipe_9596_inst 
    OutportGroup0: Block -- 
      signal data_in: std_logic_vector(143 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_d_cmd_pipe_9596_inst_req_0;
      WPIPE_d_cmd_pipe_9596_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_d_cmd_pipe_9596_inst_req_1;
      WPIPE_d_cmd_pipe_9596_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      gI: SplitGuardInterface generic map(name => "gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      data_in <= d_cmd_9595;
      d_cmd_pipe_write_0: OutputPortRevised -- 
        generic map ( name => "d_cmd_pipe", data_width => 144, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => d_cmd_pipe_pipe_write_req(0),
          oack => d_cmd_pipe_pipe_write_ack(0),
          odata => d_cmd_pipe_pipe_write_data(143 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_e_cmd_pipe_9564_inst 
    OutportGroup1: Block -- 
      signal data_in: std_logic_vector(143 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_e_cmd_pipe_9564_inst_req_0;
      WPIPE_e_cmd_pipe_9564_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_e_cmd_pipe_9564_inst_req_1;
      WPIPE_e_cmd_pipe_9564_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      gI: SplitGuardInterface generic map(name => "gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      data_in <= e_cmd_9563;
      e_cmd_pipe_write_1: OutputPortRevised -- 
        generic map ( name => "e_cmd_pipe", data_width => 144, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => e_cmd_pipe_pipe_write_req(0),
          oack => e_cmd_pipe_pipe_write_ack(0),
          odata => e_cmd_pipe_pipe_write_data(143 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared outport operator group (2) : WPIPE_status_out_9574_inst WPIPE_status_out_9542_inst 
    OutportGroup2: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal sample_req, sample_ack : BooleanArray( 1 downto 0);
      signal update_req, update_ack : BooleanArray( 1 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 1 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      sample_req_unguarded(1) <= WPIPE_status_out_9574_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_status_out_9542_inst_req_0;
      WPIPE_status_out_9574_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_status_out_9542_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(1) <= WPIPE_status_out_9574_inst_req_1;
      update_req_unguarded(0) <= WPIPE_status_out_9542_inst_req_1;
      WPIPE_status_out_9574_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_status_out_9542_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      gI: SplitGuardInterface generic map(name => "gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      data_in <= konst_9575_wire_constant & konst_9543_wire_constant;
      status_out_write_2: OutputPortRevised -- 
        generic map ( name => "status_out", data_width => 64, num_reqs => 2, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => status_out_pipe_write_req(0),
          oack => status_out_pipe_write_ack(0),
          odata => status_out_pipe_write_data(63 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 2
    -- 
  end Block; -- data_path
  -- 
end c_block_daemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library work;
use work.ahir_system_global_package.all;
entity d_block_daemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    d_cmd_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    d_cmd_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    d_cmd_pipe_pipe_read_data : in   std_logic_vector(143 downto 0);
    d_in_buf_pipe_read_req : out  std_logic_vector(0 downto 0);
    d_in_buf_pipe_read_ack : in   std_logic_vector(0 downto 0);
    d_in_buf_pipe_read_data : in   std_logic_vector(127 downto 0);
    d_block_done_pipe_write_req : out  std_logic_vector(0 downto 0);
    d_block_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
    d_block_done_pipe_write_data : out  std_logic_vector(0 downto 0);
    d_out_buf_pipe_write_req : out  std_logic_vector(0 downto 0);
    d_out_buf_pipe_write_ack : in   std_logic_vector(0 downto 0);
    d_out_buf_pipe_write_data : out  std_logic_vector(127 downto 0);
    key_expand_single_call_reqs : out  std_logic_vector(0 downto 0);
    key_expand_single_call_acks : in   std_logic_vector(0 downto 0);
    key_expand_single_call_data : out  std_logic_vector(135 downto 0);
    key_expand_single_call_tag  :  out  std_logic_vector(3 downto 0);
    key_expand_single_return_reqs : out  std_logic_vector(0 downto 0);
    key_expand_single_return_acks : in   std_logic_vector(0 downto 0);
    key_expand_single_return_data : in   std_logic_vector(135 downto 0);
    key_expand_single_return_tag :  in   std_logic_vector(3 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity d_block_daemon;
architecture d_block_daemon_arch of d_block_daemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal d_block_daemon_CP_6409_start: Boolean;
  signal d_block_daemon_CP_6409_symbol: Boolean;
  -- volatile/operator module components. 
  component key_expand_single is -- 
    generic (tag_length : integer); 
    port ( -- 
      K_in : in  std_logic_vector(127 downto 0);
      Round_C : in  std_logic_vector(7 downto 0);
      K_out : out  std_logic_vector(127 downto 0);
      nRound_C : out  std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component dec_round_Operator is -- 
    port ( -- 
      sample_req: in boolean;
      sample_ack: out boolean;
      update_req: in boolean;
      update_ack: out boolean;
      round_in : in  std_logic_vector(127 downto 0);
      key_in : in  std_logic_vector(127 downto 0);
      l_round : in  std_logic_vector(0 downto 0);
      round_out : out  std_logic_vector(127 downto 0);
      clk, reset: in std_logic
      -- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal RPIPE_d_cmd_pipe_12838_inst_ack_1 : boolean;
  signal RPIPE_d_cmd_pipe_12838_inst_req_1 : boolean;
  signal RPIPE_d_cmd_pipe_12838_inst_ack_0 : boolean;
  signal RPIPE_d_cmd_pipe_12838_inst_req_0 : boolean;
  signal WPIPE_d_block_done_12833_inst_ack_1 : boolean;
  signal WPIPE_d_block_done_12833_inst_req_1 : boolean;
  signal call_stmt_12917_call_req_0 : boolean;
  signal WPIPE_d_block_done_12833_inst_ack_0 : boolean;
  signal WPIPE_d_block_done_12833_inst_req_0 : boolean;
  signal call_stmt_12917_call_ack_0 : boolean;
  signal call_stmt_12907_call_req_0 : boolean;
  signal call_stmt_12917_call_ack_1 : boolean;
  signal call_stmt_12907_call_ack_1 : boolean;
  signal W_K9_12940_delayed_1_12942_inst_req_1 : boolean;
  signal W_K9_12940_delayed_1_12942_inst_ack_0 : boolean;
  signal W_K9_12940_delayed_1_12942_inst_req_0 : boolean;
  signal call_stmt_12907_call_ack_0 : boolean;
  signal call_stmt_12917_call_req_1 : boolean;
  signal do_while_stmt_12924_branch_req_0 : boolean;
  signal RPIPE_d_in_buf_12932_inst_ack_0 : boolean;
  signal RPIPE_d_in_buf_12932_inst_req_0 : boolean;
  signal W_K10_12936_delayed_1_12934_inst_ack_1 : boolean;
  signal W_K9_12940_delayed_1_12942_inst_ack_1 : boolean;
  signal W_K10_12936_delayed_1_12934_inst_req_1 : boolean;
  signal call_stmt_12912_call_ack_1 : boolean;
  signal call_stmt_12912_call_req_1 : boolean;
  signal if_stmt_12852_branch_req_0 : boolean;
  signal if_stmt_12852_branch_ack_1 : boolean;
  signal call_stmt_12912_call_ack_0 : boolean;
  signal if_stmt_12852_branch_ack_0 : boolean;
  signal n_count_var_13029_12929_buf_ack_1 : boolean;
  signal call_stmt_12912_call_req_0 : boolean;
  signal n_count_var_13029_12929_buf_req_1 : boolean;
  signal call_stmt_12872_call_req_0 : boolean;
  signal call_stmt_12872_call_ack_0 : boolean;
  signal call_stmt_12872_call_req_1 : boolean;
  signal call_stmt_12872_call_ack_1 : boolean;
  signal n_count_var_13029_12929_buf_ack_0 : boolean;
  signal n_count_var_13029_12929_buf_req_0 : boolean;
  signal phi_stmt_12926_ack_0 : boolean;
  signal call_stmt_12877_call_req_0 : boolean;
  signal call_stmt_12877_call_ack_0 : boolean;
  signal call_stmt_12877_call_req_1 : boolean;
  signal call_stmt_12877_call_ack_1 : boolean;
  signal W_K10_12936_delayed_1_12934_inst_ack_0 : boolean;
  signal W_K10_12936_delayed_1_12934_inst_req_0 : boolean;
  signal call_stmt_12882_call_req_0 : boolean;
  signal call_stmt_12882_call_ack_0 : boolean;
  signal call_stmt_12882_call_req_1 : boolean;
  signal call_stmt_12882_call_ack_1 : boolean;
  signal RPIPE_d_in_buf_12932_inst_ack_1 : boolean;
  signal call_stmt_12887_call_req_0 : boolean;
  signal call_stmt_12887_call_ack_0 : boolean;
  signal call_stmt_12887_call_req_1 : boolean;
  signal call_stmt_12887_call_ack_1 : boolean;
  signal phi_stmt_12926_req_0 : boolean;
  signal RPIPE_d_in_buf_12932_inst_req_1 : boolean;
  signal call_stmt_12892_call_req_0 : boolean;
  signal call_stmt_12892_call_ack_0 : boolean;
  signal call_stmt_12907_call_req_1 : boolean;
  signal call_stmt_12892_call_req_1 : boolean;
  signal call_stmt_12892_call_ack_1 : boolean;
  signal phi_stmt_12926_req_1 : boolean;
  signal call_stmt_12897_call_req_0 : boolean;
  signal call_stmt_12897_call_ack_0 : boolean;
  signal call_stmt_12897_call_req_1 : boolean;
  signal call_stmt_12897_call_ack_1 : boolean;
  signal call_stmt_12902_call_req_0 : boolean;
  signal call_stmt_12902_call_ack_0 : boolean;
  signal call_stmt_12902_call_req_1 : boolean;
  signal call_stmt_12902_call_ack_1 : boolean;
  signal call_stmt_12949_call_req_0 : boolean;
  signal call_stmt_12949_call_ack_0 : boolean;
  signal call_stmt_12949_call_req_1 : boolean;
  signal call_stmt_12949_call_ack_1 : boolean;
  signal W_K8_12945_delayed_2_12950_inst_req_0 : boolean;
  signal W_K8_12945_delayed_2_12950_inst_ack_0 : boolean;
  signal W_K8_12945_delayed_2_12950_inst_req_1 : boolean;
  signal W_K8_12945_delayed_2_12950_inst_ack_1 : boolean;
  signal call_stmt_12957_call_req_0 : boolean;
  signal call_stmt_12957_call_ack_0 : boolean;
  signal call_stmt_12957_call_req_1 : boolean;
  signal call_stmt_12957_call_ack_1 : boolean;
  signal W_K7_12950_delayed_3_12958_inst_req_0 : boolean;
  signal W_K7_12950_delayed_3_12958_inst_ack_0 : boolean;
  signal W_K7_12950_delayed_3_12958_inst_req_1 : boolean;
  signal W_K7_12950_delayed_3_12958_inst_ack_1 : boolean;
  signal call_stmt_12965_call_req_0 : boolean;
  signal call_stmt_12965_call_ack_0 : boolean;
  signal call_stmt_12965_call_req_1 : boolean;
  signal call_stmt_12965_call_ack_1 : boolean;
  signal W_K6_12955_delayed_4_12966_inst_req_0 : boolean;
  signal W_K6_12955_delayed_4_12966_inst_ack_0 : boolean;
  signal W_K6_12955_delayed_4_12966_inst_req_1 : boolean;
  signal W_K6_12955_delayed_4_12966_inst_ack_1 : boolean;
  signal call_stmt_12973_call_req_0 : boolean;
  signal call_stmt_12973_call_ack_0 : boolean;
  signal call_stmt_12973_call_req_1 : boolean;
  signal call_stmt_12973_call_ack_1 : boolean;
  signal W_K5_12960_delayed_5_12974_inst_req_0 : boolean;
  signal W_K5_12960_delayed_5_12974_inst_ack_0 : boolean;
  signal W_K5_12960_delayed_5_12974_inst_req_1 : boolean;
  signal W_K5_12960_delayed_5_12974_inst_ack_1 : boolean;
  signal call_stmt_12981_call_req_0 : boolean;
  signal call_stmt_12981_call_ack_0 : boolean;
  signal call_stmt_12981_call_req_1 : boolean;
  signal call_stmt_12981_call_ack_1 : boolean;
  signal W_K4_12965_delayed_6_12982_inst_req_0 : boolean;
  signal W_K4_12965_delayed_6_12982_inst_ack_0 : boolean;
  signal W_K4_12965_delayed_6_12982_inst_req_1 : boolean;
  signal W_K4_12965_delayed_6_12982_inst_ack_1 : boolean;
  signal call_stmt_12989_call_req_0 : boolean;
  signal call_stmt_12989_call_ack_0 : boolean;
  signal call_stmt_12989_call_req_1 : boolean;
  signal call_stmt_12989_call_ack_1 : boolean;
  signal phi_stmt_12919_req_0 : boolean;
  signal W_K3_12970_delayed_7_12990_inst_req_0 : boolean;
  signal W_K3_12970_delayed_7_12990_inst_ack_0 : boolean;
  signal W_K3_12970_delayed_7_12990_inst_req_1 : boolean;
  signal W_K3_12970_delayed_7_12990_inst_ack_1 : boolean;
  signal d_new_count_13047_12922_buf_req_0 : boolean;
  signal d_new_count_13047_12922_buf_ack_0 : boolean;
  signal d_new_count_13047_12922_buf_req_1 : boolean;
  signal phi_stmt_12859_req_0 : boolean;
  signal countA_12863_12921_buf_req_1 : boolean;
  signal countA_12863_12921_buf_ack_1 : boolean;
  signal phi_stmt_12863_req_1 : boolean;
  signal call_stmt_12997_call_req_0 : boolean;
  signal call_stmt_12997_call_ack_0 : boolean;
  signal call_stmt_12997_call_req_1 : boolean;
  signal call_stmt_12997_call_ack_1 : boolean;
  signal d_init_key_12851_12861_buf_ack_1 : boolean;
  signal countA_12863_12921_buf_req_0 : boolean;
  signal countA_12863_12921_buf_ack_0 : boolean;
  signal d_init_key_12851_12861_buf_req_1 : boolean;
  signal W_K2_12975_delayed_8_12998_inst_req_0 : boolean;
  signal W_K2_12975_delayed_8_12998_inst_ack_0 : boolean;
  signal W_K2_12975_delayed_8_12998_inst_req_1 : boolean;
  signal W_K2_12975_delayed_8_12998_inst_ack_1 : boolean;
  signal d_init_key_12851_12861_buf_ack_0 : boolean;
  signal d_new_count_13047_12866_buf_ack_1 : boolean;
  signal phi_stmt_12863_req_0 : boolean;
  signal call_stmt_13005_call_req_0 : boolean;
  signal call_stmt_13005_call_ack_0 : boolean;
  signal call_stmt_13005_call_req_1 : boolean;
  signal call_stmt_13005_call_ack_1 : boolean;
  signal d_init_key_12851_12861_buf_req_0 : boolean;
  signal d_init_count_12847_12865_buf_ack_1 : boolean;
  signal d_init_count_12847_12865_buf_req_1 : boolean;
  signal W_K1_12980_delayed_9_13006_inst_req_0 : boolean;
  signal W_K1_12980_delayed_9_13006_inst_ack_0 : boolean;
  signal W_K1_12980_delayed_9_13006_inst_req_1 : boolean;
  signal W_K1_12980_delayed_9_13006_inst_ack_1 : boolean;
  signal d_new_count_13047_12922_buf_ack_1 : boolean;
  signal phi_stmt_12919_req_1 : boolean;
  signal phi_stmt_12863_ack_0 : boolean;
  signal d_new_count_13047_12866_buf_req_1 : boolean;
  signal d_init_count_12847_12865_buf_ack_0 : boolean;
  signal d_init_count_12847_12865_buf_req_0 : boolean;
  signal phi_stmt_12859_req_1 : boolean;
  signal d_new_key_13051_12862_buf_ack_1 : boolean;
  signal d_new_key_13051_12862_buf_req_1 : boolean;
  signal call_stmt_13013_call_req_0 : boolean;
  signal call_stmt_13013_call_ack_0 : boolean;
  signal call_stmt_13013_call_req_1 : boolean;
  signal call_stmt_13013_call_ack_1 : boolean;
  signal W_K0_12985_delayed_10_13014_inst_req_0 : boolean;
  signal W_K0_12985_delayed_10_13014_inst_ack_0 : boolean;
  signal W_K0_12985_delayed_10_13014_inst_req_1 : boolean;
  signal W_K0_12985_delayed_10_13014_inst_ack_1 : boolean;
  signal phi_stmt_12859_ack_0 : boolean;
  signal d_new_key_13051_12862_buf_ack_0 : boolean;
  signal d_new_count_13047_12866_buf_ack_0 : boolean;
  signal d_new_count_13047_12866_buf_req_0 : boolean;
  signal call_stmt_13021_call_req_0 : boolean;
  signal call_stmt_13021_call_ack_0 : boolean;
  signal call_stmt_13021_call_req_1 : boolean;
  signal call_stmt_13021_call_ack_1 : boolean;
  signal if_stmt_13052_branch_ack_0 : boolean;
  signal if_stmt_13052_branch_ack_1 : boolean;
  signal WPIPE_d_out_buf_13022_inst_req_0 : boolean;
  signal WPIPE_d_out_buf_13022_inst_ack_0 : boolean;
  signal WPIPE_d_out_buf_13022_inst_req_1 : boolean;
  signal WPIPE_d_out_buf_13022_inst_ack_1 : boolean;
  signal d_new_key_13051_12862_buf_req_0 : boolean;
  signal if_stmt_13052_branch_req_0 : boolean;
  signal ADD_u15_u15_13028_inst_req_0 : boolean;
  signal ADD_u15_u15_13028_inst_ack_0 : boolean;
  signal ADD_u15_u15_13028_inst_req_1 : boolean;
  signal ADD_u15_u15_13028_inst_ack_1 : boolean;
  signal do_while_stmt_12924_branch_ack_0 : boolean;
  signal do_while_stmt_12924_branch_ack_1 : boolean;
  signal WPIPE_d_block_done_13034_inst_req_0 : boolean;
  signal WPIPE_d_block_done_13034_inst_ack_0 : boolean;
  signal WPIPE_d_block_done_13034_inst_req_1 : boolean;
  signal WPIPE_d_block_done_13034_inst_ack_1 : boolean;
  signal RPIPE_d_cmd_pipe_13038_inst_req_0 : boolean;
  signal RPIPE_d_cmd_pipe_13038_inst_ack_0 : boolean;
  signal RPIPE_d_cmd_pipe_13038_inst_req_1 : boolean;
  signal RPIPE_d_cmd_pipe_13038_inst_ack_1 : boolean;
  signal phi_stmt_12919_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "d_block_daemon_input_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      bypass_flag => true,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  d_block_daemon_CP_6409_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "d_block_daemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= d_block_daemon_CP_6409_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= d_block_daemon_CP_6409_start & tag_ilock_write_ack_symbol;
    gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= d_block_daemon_CP_6409_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  d_block_daemon_CP_6409: Block -- control-path 
    signal d_block_daemon_CP_6409_elements: BooleanArray(249 downto 0);
    -- 
  begin -- 
    d_block_daemon_CP_6409_elements(0) <= d_block_daemon_CP_6409_start;
    -- unreachable exit of control-path
    d_block_daemon_CP_6409_symbol <= false;
    -- CP-element group 0:  transition  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (2) 
      -- CP-element group 0: 	 branch_block_stmt_12832/$entry
      -- CP-element group 0: 	 $entry
      -- 
    -- CP-element group 1:  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	14 
    -- CP-element group 1:  members (2) 
      -- CP-element group 1: 	 branch_block_stmt_12832/assign_stmt_12835__entry__
      -- CP-element group 1: 	 branch_block_stmt_12832/branch_block_stmt_12832__entry__
      -- 
    d_block_daemon_CP_6409_elements(1) <= d_block_daemon_CP_6409_elements(0);
    -- CP-element group 2:  branch  place  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	16 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	210 
    -- CP-element group 2: 	211 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_12832/merge_stmt_12836__entry__
      -- CP-element group 2: 	 branch_block_stmt_12832/assign_stmt_12835__exit__
      -- 
    d_block_daemon_CP_6409_elements(2) <= d_block_daemon_CP_6409_elements(16);
    -- CP-element group 3:  merge  place  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	214 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	17 
    -- CP-element group 3:  members (2) 
      -- CP-element group 3: 	 branch_block_stmt_12832/assign_stmt_12839__entry__
      -- CP-element group 3: 	 branch_block_stmt_12832/merge_stmt_12836__exit__
      -- 
    d_block_daemon_CP_6409_elements(3) <= d_block_daemon_CP_6409_elements(214);
    -- CP-element group 4:  place  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	19 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	20 
    -- CP-element group 4:  members (2) 
      -- CP-element group 4: 	 branch_block_stmt_12832/assign_stmt_12843_to_assign_stmt_12851__entry__
      -- CP-element group 4: 	 branch_block_stmt_12832/assign_stmt_12839__exit__
      -- 
    d_block_daemon_CP_6409_elements(4) <= d_block_daemon_CP_6409_elements(19);
    -- CP-element group 5:  branch  place  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	20 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	21 
    -- CP-element group 5: 	22 
    -- CP-element group 5:  members (2) 
      -- CP-element group 5: 	 branch_block_stmt_12832/if_stmt_12852__entry__
      -- CP-element group 5: 	 branch_block_stmt_12832/assign_stmt_12843_to_assign_stmt_12851__exit__
      -- 
    d_block_daemon_CP_6409_elements(5) <= d_block_daemon_CP_6409_elements(20);
    -- CP-element group 6:  merge  branch  place  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	27 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	215 
    -- CP-element group 6: 	216 
    -- CP-element group 6:  members (2) 
      -- CP-element group 6: 	 branch_block_stmt_12832/merge_stmt_12858__entry__
      -- CP-element group 6: 	 branch_block_stmt_12832/if_stmt_12852__exit__
      -- 
    d_block_daemon_CP_6409_elements(6) <= d_block_daemon_CP_6409_elements(27);
    -- CP-element group 7:  merge  place  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	236 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	29 
    -- CP-element group 7:  members (2) 
      -- CP-element group 7: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917__entry__
      -- CP-element group 7: 	 branch_block_stmt_12832/merge_stmt_12858__exit__
      -- 
    d_block_daemon_CP_6409_elements(7) <= d_block_daemon_CP_6409_elements(236);
    -- CP-element group 8:  branch  place  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	49 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	237 
    -- CP-element group 8: 	238 
    -- CP-element group 8:  members (2) 
      -- CP-element group 8: 	 branch_block_stmt_12832/merge_stmt_12918__entry__
      -- CP-element group 8: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917__exit__
      -- 
    d_block_daemon_CP_6409_elements(8) <= d_block_daemon_CP_6409_elements(49);
    -- CP-element group 9:  merge  place  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	248 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	50 
    -- CP-element group 9:  members (2) 
      -- CP-element group 9: 	 branch_block_stmt_12832/do_while_stmt_12924__entry__
      -- CP-element group 9: 	 branch_block_stmt_12832/merge_stmt_12918__exit__
      -- 
    d_block_daemon_CP_6409_elements(9) <= d_block_daemon_CP_6409_elements(248);
    -- CP-element group 10:  place  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	193 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	194 
    -- CP-element group 10:  members (2) 
      -- CP-element group 10: 	 branch_block_stmt_12832/assign_stmt_13036__entry__
      -- CP-element group 10: 	 branch_block_stmt_12832/do_while_stmt_12924__exit__
      -- 
    d_block_daemon_CP_6409_elements(10) <= d_block_daemon_CP_6409_elements(193);
    -- CP-element group 11:  place  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	196 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	197 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_12832/assign_stmt_13039__entry__
      -- CP-element group 11: 	 branch_block_stmt_12832/assign_stmt_13036__exit__
      -- 
    d_block_daemon_CP_6409_elements(11) <= d_block_daemon_CP_6409_elements(196);
    -- CP-element group 12:  place  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	199 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	200 
    -- CP-element group 12:  members (2) 
      -- CP-element group 12: 	 branch_block_stmt_12832/assign_stmt_13043_to_assign_stmt_13051__entry__
      -- CP-element group 12: 	 branch_block_stmt_12832/assign_stmt_13039__exit__
      -- 
    d_block_daemon_CP_6409_elements(12) <= d_block_daemon_CP_6409_elements(199);
    -- CP-element group 13:  branch  place  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	200 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	201 
    -- CP-element group 13: 	202 
    -- CP-element group 13:  members (2) 
      -- CP-element group 13: 	 branch_block_stmt_12832/if_stmt_13052__entry__
      -- CP-element group 13: 	 branch_block_stmt_12832/assign_stmt_13043_to_assign_stmt_13051__exit__
      -- 
    d_block_daemon_CP_6409_elements(13) <= d_block_daemon_CP_6409_elements(200);
    -- CP-element group 14:  transition  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	1 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (4) 
      -- CP-element group 14: 	 branch_block_stmt_12832/assign_stmt_12835/WPIPE_d_block_done_12833_Sample/req
      -- CP-element group 14: 	 branch_block_stmt_12832/assign_stmt_12835/WPIPE_d_block_done_12833_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_12832/assign_stmt_12835/WPIPE_d_block_done_12833_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_12832/assign_stmt_12835/$entry
      -- 
    req_6453_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6453_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_6409_elements(14), ack => WPIPE_d_block_done_12833_inst_req_0); -- 
    d_block_daemon_CP_6409_elements(14) <= d_block_daemon_CP_6409_elements(1);
    -- CP-element group 15:  transition  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (6) 
      -- CP-element group 15: 	 branch_block_stmt_12832/assign_stmt_12835/WPIPE_d_block_done_12833_Update/req
      -- CP-element group 15: 	 branch_block_stmt_12832/assign_stmt_12835/WPIPE_d_block_done_12833_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_12832/assign_stmt_12835/WPIPE_d_block_done_12833_Sample/ack
      -- CP-element group 15: 	 branch_block_stmt_12832/assign_stmt_12835/WPIPE_d_block_done_12833_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_12832/assign_stmt_12835/WPIPE_d_block_done_12833_update_start_
      -- CP-element group 15: 	 branch_block_stmt_12832/assign_stmt_12835/WPIPE_d_block_done_12833_sample_completed_
      -- 
    ack_6454_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_d_block_done_12833_inst_ack_0, ack => d_block_daemon_CP_6409_elements(15)); -- 
    req_6458_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6458_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_6409_elements(15), ack => WPIPE_d_block_done_12833_inst_req_1); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	2 
    -- CP-element group 16:  members (4) 
      -- CP-element group 16: 	 branch_block_stmt_12832/assign_stmt_12835/WPIPE_d_block_done_12833_Update/ack
      -- CP-element group 16: 	 branch_block_stmt_12832/assign_stmt_12835/WPIPE_d_block_done_12833_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_12832/assign_stmt_12835/WPIPE_d_block_done_12833_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_12832/assign_stmt_12835/$exit
      -- 
    ack_6459_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_d_block_done_12833_inst_ack_1, ack => d_block_daemon_CP_6409_elements(16)); -- 
    -- CP-element group 17:  transition  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	3 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (4) 
      -- CP-element group 17: 	 branch_block_stmt_12832/assign_stmt_12839/RPIPE_d_cmd_pipe_12838_Sample/rr
      -- CP-element group 17: 	 branch_block_stmt_12832/assign_stmt_12839/RPIPE_d_cmd_pipe_12838_Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_12832/assign_stmt_12839/RPIPE_d_cmd_pipe_12838_sample_start_
      -- CP-element group 17: 	 branch_block_stmt_12832/assign_stmt_12839/$entry
      -- 
    rr_6470_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6470_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_6409_elements(17), ack => RPIPE_d_cmd_pipe_12838_inst_req_0); -- 
    d_block_daemon_CP_6409_elements(17) <= d_block_daemon_CP_6409_elements(3);
    -- CP-element group 18:  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (6) 
      -- CP-element group 18: 	 branch_block_stmt_12832/assign_stmt_12839/RPIPE_d_cmd_pipe_12838_Update/cr
      -- CP-element group 18: 	 branch_block_stmt_12832/assign_stmt_12839/RPIPE_d_cmd_pipe_12838_Update/$entry
      -- CP-element group 18: 	 branch_block_stmt_12832/assign_stmt_12839/RPIPE_d_cmd_pipe_12838_Sample/ra
      -- CP-element group 18: 	 branch_block_stmt_12832/assign_stmt_12839/RPIPE_d_cmd_pipe_12838_Sample/$exit
      -- CP-element group 18: 	 branch_block_stmt_12832/assign_stmt_12839/RPIPE_d_cmd_pipe_12838_update_start_
      -- CP-element group 18: 	 branch_block_stmt_12832/assign_stmt_12839/RPIPE_d_cmd_pipe_12838_sample_completed_
      -- 
    ra_6471_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_d_cmd_pipe_12838_inst_ack_0, ack => d_block_daemon_CP_6409_elements(18)); -- 
    cr_6475_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6475_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_6409_elements(18), ack => RPIPE_d_cmd_pipe_12838_inst_req_1); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	4 
    -- CP-element group 19:  members (4) 
      -- CP-element group 19: 	 branch_block_stmt_12832/assign_stmt_12839/RPIPE_d_cmd_pipe_12838_Update/ca
      -- CP-element group 19: 	 branch_block_stmt_12832/assign_stmt_12839/RPIPE_d_cmd_pipe_12838_Update/$exit
      -- CP-element group 19: 	 branch_block_stmt_12832/assign_stmt_12839/RPIPE_d_cmd_pipe_12838_update_completed_
      -- CP-element group 19: 	 branch_block_stmt_12832/assign_stmt_12839/$exit
      -- 
    ca_6476_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_d_cmd_pipe_12838_inst_ack_1, ack => d_block_daemon_CP_6409_elements(19)); -- 
    -- CP-element group 20:  join  fork  transition  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	4 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	5 
    -- CP-element group 20:  members (50) 
      -- CP-element group 20: 	 branch_block_stmt_12832/assign_stmt_12843_to_assign_stmt_12851/$exit
      -- CP-element group 20: 	 branch_block_stmt_12832/assign_stmt_12843_to_assign_stmt_12851/$entry
      -- CP-element group 20: 	 branch_block_stmt_12832/assign_stmt_12843_to_assign_stmt_12851/slice_12842_sample_start_
      -- CP-element group 20: 	 branch_block_stmt_12832/assign_stmt_12843_to_assign_stmt_12851/slice_12842_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_12832/assign_stmt_12843_to_assign_stmt_12851/slice_12842_update_start_
      -- CP-element group 20: 	 branch_block_stmt_12832/assign_stmt_12843_to_assign_stmt_12851/slice_12842_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_12832/assign_stmt_12843_to_assign_stmt_12851/R_d_init_cmd_12841_sample_start_
      -- CP-element group 20: 	 branch_block_stmt_12832/assign_stmt_12843_to_assign_stmt_12851/R_d_init_cmd_12841_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_12832/assign_stmt_12843_to_assign_stmt_12851/R_d_init_cmd_12841_update_start_
      -- CP-element group 20: 	 branch_block_stmt_12832/assign_stmt_12843_to_assign_stmt_12851/R_d_init_cmd_12841_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_12832/assign_stmt_12843_to_assign_stmt_12851/slice_12842_Sample/$entry
      -- CP-element group 20: 	 branch_block_stmt_12832/assign_stmt_12843_to_assign_stmt_12851/slice_12842_Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_12832/assign_stmt_12843_to_assign_stmt_12851/slice_12842_Sample/rr
      -- CP-element group 20: 	 branch_block_stmt_12832/assign_stmt_12843_to_assign_stmt_12851/slice_12842_Sample/ra
      -- CP-element group 20: 	 branch_block_stmt_12832/assign_stmt_12843_to_assign_stmt_12851/slice_12842_Update/$entry
      -- CP-element group 20: 	 branch_block_stmt_12832/assign_stmt_12843_to_assign_stmt_12851/slice_12842_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_12832/assign_stmt_12843_to_assign_stmt_12851/slice_12842_Update/cr
      -- CP-element group 20: 	 branch_block_stmt_12832/assign_stmt_12843_to_assign_stmt_12851/slice_12842_Update/ca
      -- CP-element group 20: 	 branch_block_stmt_12832/assign_stmt_12843_to_assign_stmt_12851/slice_12846_sample_start_
      -- CP-element group 20: 	 branch_block_stmt_12832/assign_stmt_12843_to_assign_stmt_12851/slice_12846_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_12832/assign_stmt_12843_to_assign_stmt_12851/slice_12846_update_start_
      -- CP-element group 20: 	 branch_block_stmt_12832/assign_stmt_12843_to_assign_stmt_12851/slice_12846_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_12832/assign_stmt_12843_to_assign_stmt_12851/R_d_init_cmd_12845_sample_start_
      -- CP-element group 20: 	 branch_block_stmt_12832/assign_stmt_12843_to_assign_stmt_12851/R_d_init_cmd_12845_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_12832/assign_stmt_12843_to_assign_stmt_12851/R_d_init_cmd_12845_update_start_
      -- CP-element group 20: 	 branch_block_stmt_12832/assign_stmt_12843_to_assign_stmt_12851/R_d_init_cmd_12845_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_12832/assign_stmt_12843_to_assign_stmt_12851/slice_12846_Sample/$entry
      -- CP-element group 20: 	 branch_block_stmt_12832/assign_stmt_12843_to_assign_stmt_12851/slice_12846_Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_12832/assign_stmt_12843_to_assign_stmt_12851/slice_12846_Sample/rr
      -- CP-element group 20: 	 branch_block_stmt_12832/assign_stmt_12843_to_assign_stmt_12851/slice_12846_Sample/ra
      -- CP-element group 20: 	 branch_block_stmt_12832/assign_stmt_12843_to_assign_stmt_12851/slice_12846_Update/$entry
      -- CP-element group 20: 	 branch_block_stmt_12832/assign_stmt_12843_to_assign_stmt_12851/slice_12846_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_12832/assign_stmt_12843_to_assign_stmt_12851/slice_12846_Update/cr
      -- CP-element group 20: 	 branch_block_stmt_12832/assign_stmt_12843_to_assign_stmt_12851/slice_12846_Update/ca
      -- CP-element group 20: 	 branch_block_stmt_12832/assign_stmt_12843_to_assign_stmt_12851/slice_12850_sample_start_
      -- CP-element group 20: 	 branch_block_stmt_12832/assign_stmt_12843_to_assign_stmt_12851/slice_12850_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_12832/assign_stmt_12843_to_assign_stmt_12851/slice_12850_update_start_
      -- CP-element group 20: 	 branch_block_stmt_12832/assign_stmt_12843_to_assign_stmt_12851/slice_12850_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_12832/assign_stmt_12843_to_assign_stmt_12851/R_d_init_cmd_12849_sample_start_
      -- CP-element group 20: 	 branch_block_stmt_12832/assign_stmt_12843_to_assign_stmt_12851/R_d_init_cmd_12849_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_12832/assign_stmt_12843_to_assign_stmt_12851/R_d_init_cmd_12849_update_start_
      -- CP-element group 20: 	 branch_block_stmt_12832/assign_stmt_12843_to_assign_stmt_12851/R_d_init_cmd_12849_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_12832/assign_stmt_12843_to_assign_stmt_12851/slice_12850_Sample/$entry
      -- CP-element group 20: 	 branch_block_stmt_12832/assign_stmt_12843_to_assign_stmt_12851/slice_12850_Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_12832/assign_stmt_12843_to_assign_stmt_12851/slice_12850_Sample/rr
      -- CP-element group 20: 	 branch_block_stmt_12832/assign_stmt_12843_to_assign_stmt_12851/slice_12850_Sample/ra
      -- CP-element group 20: 	 branch_block_stmt_12832/assign_stmt_12843_to_assign_stmt_12851/slice_12850_Update/$entry
      -- CP-element group 20: 	 branch_block_stmt_12832/assign_stmt_12843_to_assign_stmt_12851/slice_12850_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_12832/assign_stmt_12843_to_assign_stmt_12851/slice_12850_Update/cr
      -- CP-element group 20: 	 branch_block_stmt_12832/assign_stmt_12843_to_assign_stmt_12851/slice_12850_Update/ca
      -- 
    d_block_daemon_CP_6409_elements(20) <= d_block_daemon_CP_6409_elements(4);
    -- CP-element group 21:  transition  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	5 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_12832/if_stmt_12852_dead_link/$entry
      -- 
    d_block_daemon_CP_6409_elements(21) <= d_block_daemon_CP_6409_elements(5);
    -- CP-element group 22:  transition  output  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	5 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	23 
    -- CP-element group 22:  members (17) 
      -- CP-element group 22: 	 branch_block_stmt_12832/if_stmt_12852_eval_test/$entry
      -- CP-element group 22: 	 branch_block_stmt_12832/if_stmt_12852_eval_test/$exit
      -- CP-element group 22: 	 branch_block_stmt_12832/if_stmt_12852_eval_test/EQ_u1_u1_12855/$entry
      -- CP-element group 22: 	 branch_block_stmt_12832/if_stmt_12852_eval_test/EQ_u1_u1_12855/$exit
      -- CP-element group 22: 	 branch_block_stmt_12832/if_stmt_12852_eval_test/EQ_u1_u1_12855/EQ_u1_u1_12855_inputs/$entry
      -- CP-element group 22: 	 branch_block_stmt_12832/if_stmt_12852_eval_test/EQ_u1_u1_12855/EQ_u1_u1_12855_inputs/$exit
      -- CP-element group 22: 	 branch_block_stmt_12832/if_stmt_12852_eval_test/EQ_u1_u1_12855/SplitProtocol/$entry
      -- CP-element group 22: 	 branch_block_stmt_12832/if_stmt_12852_eval_test/EQ_u1_u1_12855/SplitProtocol/$exit
      -- CP-element group 22: 	 branch_block_stmt_12832/if_stmt_12852_eval_test/EQ_u1_u1_12855/SplitProtocol/Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_12832/if_stmt_12852_eval_test/EQ_u1_u1_12855/SplitProtocol/Sample/$exit
      -- CP-element group 22: 	 branch_block_stmt_12832/if_stmt_12852_eval_test/EQ_u1_u1_12855/SplitProtocol/Sample/rr
      -- CP-element group 22: 	 branch_block_stmt_12832/if_stmt_12852_eval_test/EQ_u1_u1_12855/SplitProtocol/Sample/ra
      -- CP-element group 22: 	 branch_block_stmt_12832/if_stmt_12852_eval_test/EQ_u1_u1_12855/SplitProtocol/Update/$entry
      -- CP-element group 22: 	 branch_block_stmt_12832/if_stmt_12852_eval_test/EQ_u1_u1_12855/SplitProtocol/Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_12832/if_stmt_12852_eval_test/EQ_u1_u1_12855/SplitProtocol/Update/cr
      -- CP-element group 22: 	 branch_block_stmt_12832/if_stmt_12852_eval_test/EQ_u1_u1_12855/SplitProtocol/Update/ca
      -- CP-element group 22: 	 branch_block_stmt_12832/if_stmt_12852_eval_test/branch_req
      -- 
    branch_req_6560_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_6560_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_6409_elements(22), ack => if_stmt_12852_branch_req_0); -- 
    d_block_daemon_CP_6409_elements(22) <= d_block_daemon_CP_6409_elements(5);
    -- CP-element group 23:  branch  place  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	22 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	24 
    -- CP-element group 23: 	26 
    -- CP-element group 23:  members (1) 
      -- CP-element group 23: 	 branch_block_stmt_12832/EQ_u1_u1_12855_place
      -- 
    d_block_daemon_CP_6409_elements(23) <= d_block_daemon_CP_6409_elements(22);
    -- CP-element group 24:  transition  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	23 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24:  members (1) 
      -- CP-element group 24: 	 branch_block_stmt_12832/if_stmt_12852_if_link/$entry
      -- 
    d_block_daemon_CP_6409_elements(24) <= d_block_daemon_CP_6409_elements(23);
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	24 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	28 
    -- CP-element group 25:  members (2) 
      -- CP-element group 25: 	 branch_block_stmt_12832/if_stmt_12852_if_link/$exit
      -- CP-element group 25: 	 branch_block_stmt_12832/if_stmt_12852_if_link/if_choice_transition
      -- 
    if_choice_transition_6565_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_12852_branch_ack_1, ack => d_block_daemon_CP_6409_elements(25)); -- 
    -- CP-element group 26:  transition  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	23 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	27 
    -- CP-element group 26:  members (1) 
      -- CP-element group 26: 	 branch_block_stmt_12832/if_stmt_12852_else_link/$entry
      -- 
    d_block_daemon_CP_6409_elements(26) <= d_block_daemon_CP_6409_elements(23);
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	26 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	6 
    -- CP-element group 27:  members (2) 
      -- CP-element group 27: 	 branch_block_stmt_12832/if_stmt_12852_else_link/$exit
      -- CP-element group 27: 	 branch_block_stmt_12832/if_stmt_12852_else_link/else_choice_transition
      -- 
    else_choice_transition_6569_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_12852_branch_ack_0, ack => d_block_daemon_CP_6409_elements(27)); -- 
    -- CP-element group 28:  place  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	25 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	212 
    -- CP-element group 28:  members (1) 
      -- CP-element group 28: 	 branch_block_stmt_12832/NotGotCmd
      -- 
    d_block_daemon_CP_6409_elements(28) <= d_block_daemon_CP_6409_elements(25);
    -- CP-element group 29:  fork  transition  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	7 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29: 	31 
    -- CP-element group 29: 	41 
    -- CP-element group 29: 	33 
    -- CP-element group 29: 	43 
    -- CP-element group 29: 	35 
    -- CP-element group 29: 	37 
    -- CP-element group 29: 	45 
    -- CP-element group 29: 	49 
    -- CP-element group 29: 	39 
    -- CP-element group 29: 	47 
    -- CP-element group 29:  members (38) 
      -- CP-element group 29: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12917_Update/$entry
      -- CP-element group 29: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12917_Update/ccr
      -- CP-element group 29: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12912_update_start_
      -- CP-element group 29: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12917_update_start_
      -- CP-element group 29: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12907_Update/$entry
      -- CP-element group 29: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12912_Update/ccr
      -- CP-element group 29: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12912_Update/$entry
      -- CP-element group 29: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/$entry
      -- CP-element group 29: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12872_sample_start_
      -- CP-element group 29: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12872_update_start_
      -- CP-element group 29: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/R_K0_12868_sample_start_
      -- CP-element group 29: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/R_K0_12868_sample_completed_
      -- CP-element group 29: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/R_K0_12868_update_start_
      -- CP-element group 29: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/R_K0_12868_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12872_Sample/$entry
      -- CP-element group 29: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12872_Sample/crr
      -- CP-element group 29: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12872_Update/$entry
      -- CP-element group 29: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12872_Update/ccr
      -- CP-element group 29: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12877_update_start_
      -- CP-element group 29: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12877_Update/$entry
      -- CP-element group 29: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12877_Update/ccr
      -- CP-element group 29: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12882_update_start_
      -- CP-element group 29: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12882_Update/$entry
      -- CP-element group 29: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12882_Update/ccr
      -- CP-element group 29: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12887_update_start_
      -- CP-element group 29: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12887_Update/$entry
      -- CP-element group 29: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12887_Update/ccr
      -- CP-element group 29: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12892_update_start_
      -- CP-element group 29: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12892_Update/$entry
      -- CP-element group 29: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12907_Update/ccr
      -- CP-element group 29: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12892_Update/ccr
      -- CP-element group 29: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12897_update_start_
      -- CP-element group 29: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12897_Update/$entry
      -- CP-element group 29: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12897_Update/ccr
      -- CP-element group 29: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12902_update_start_
      -- CP-element group 29: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12902_Update/$entry
      -- CP-element group 29: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12902_Update/ccr
      -- CP-element group 29: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12907_update_start_
      -- 
    ccr_6590_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_6590_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_6409_elements(29), ack => call_stmt_12872_call_req_1); -- 
    crr_6585_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_6585_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_6409_elements(29), ack => call_stmt_12872_call_req_0); -- 
    ccr_6722_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_6722_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_6409_elements(29), ack => call_stmt_12902_call_req_1); -- 
    ccr_6612_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_6612_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_6409_elements(29), ack => call_stmt_12877_call_req_1); -- 
    ccr_6634_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_6634_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_6409_elements(29), ack => call_stmt_12882_call_req_1); -- 
    ccr_6656_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_6656_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_6409_elements(29), ack => call_stmt_12887_call_req_1); -- 
    ccr_6744_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_6744_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_6409_elements(29), ack => call_stmt_12907_call_req_1); -- 
    ccr_6766_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_6766_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_6409_elements(29), ack => call_stmt_12912_call_req_1); -- 
    ccr_6678_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_6678_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_6409_elements(29), ack => call_stmt_12892_call_req_1); -- 
    ccr_6700_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_6700_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_6409_elements(29), ack => call_stmt_12897_call_req_1); -- 
    ccr_6788_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_6788_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_6409_elements(29), ack => call_stmt_12917_call_req_1); -- 
    d_block_daemon_CP_6409_elements(29) <= d_block_daemon_CP_6409_elements(7);
    -- CP-element group 30:  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12872_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12872_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12872_Sample/cra
      -- 
    cra_6586_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_12872_call_ack_0, ack => d_block_daemon_CP_6409_elements(30)); -- 
    -- CP-element group 31:  join  fork  transition  input  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	29 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31:  members (14) 
      -- CP-element group 31: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12872_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12872_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12872_Update/cca
      -- CP-element group 31: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12877_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/R_K1_12873_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/R_K1_12873_sample_completed_
      -- CP-element group 31: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/R_K1_12873_update_start_
      -- CP-element group 31: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/R_K1_12873_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/R_RConstant_2_12874_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/R_RConstant_2_12874_sample_completed_
      -- CP-element group 31: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/R_RConstant_2_12874_update_start_
      -- CP-element group 31: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/R_RConstant_2_12874_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12877_Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12877_Sample/crr
      -- 
    cca_6591_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_12872_call_ack_1, ack => d_block_daemon_CP_6409_elements(31)); -- 
    crr_6607_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_6607_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_6409_elements(31), ack => call_stmt_12877_call_req_0); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12877_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12877_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12877_Sample/cra
      -- 
    cra_6608_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_12877_call_ack_0, ack => d_block_daemon_CP_6409_elements(32)); -- 
    -- CP-element group 33:  join  fork  transition  input  output  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	29 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (14) 
      -- CP-element group 33: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12877_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12877_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12877_Update/cca
      -- CP-element group 33: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12882_sample_start_
      -- CP-element group 33: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/R_K2_12878_sample_start_
      -- CP-element group 33: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/R_K2_12878_sample_completed_
      -- CP-element group 33: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/R_K2_12878_update_start_
      -- CP-element group 33: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/R_K2_12878_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/R_RConstant_3_12879_sample_start_
      -- CP-element group 33: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/R_RConstant_3_12879_sample_completed_
      -- CP-element group 33: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/R_RConstant_3_12879_update_start_
      -- CP-element group 33: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/R_RConstant_3_12879_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12882_Sample/$entry
      -- CP-element group 33: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12882_Sample/crr
      -- 
    cca_6613_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_12877_call_ack_1, ack => d_block_daemon_CP_6409_elements(33)); -- 
    crr_6629_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_6629_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_6409_elements(33), ack => call_stmt_12882_call_req_0); -- 
    -- CP-element group 34:  transition  input  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12882_sample_completed_
      -- CP-element group 34: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12882_Sample/$exit
      -- CP-element group 34: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12882_Sample/cra
      -- 
    cra_6630_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_12882_call_ack_0, ack => d_block_daemon_CP_6409_elements(34)); -- 
    -- CP-element group 35:  join  fork  transition  input  output  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	29 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	36 
    -- CP-element group 35:  members (14) 
      -- CP-element group 35: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12882_update_completed_
      -- CP-element group 35: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12882_Update/$exit
      -- CP-element group 35: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12882_Update/cca
      -- CP-element group 35: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12887_sample_start_
      -- CP-element group 35: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/R_K3_12883_sample_start_
      -- CP-element group 35: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/R_K3_12883_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/R_K3_12883_update_start_
      -- CP-element group 35: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/R_K3_12883_update_completed_
      -- CP-element group 35: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/R_RConstant_4_12884_sample_start_
      -- CP-element group 35: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/R_RConstant_4_12884_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/R_RConstant_4_12884_update_start_
      -- CP-element group 35: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/R_RConstant_4_12884_update_completed_
      -- CP-element group 35: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12887_Sample/$entry
      -- CP-element group 35: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12887_Sample/crr
      -- 
    cca_6635_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_12882_call_ack_1, ack => d_block_daemon_CP_6409_elements(35)); -- 
    crr_6651_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_6651_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_6409_elements(35), ack => call_stmt_12887_call_req_0); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	35 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12887_sample_completed_
      -- CP-element group 36: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12887_Sample/$exit
      -- CP-element group 36: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12887_Sample/cra
      -- 
    cra_6652_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_12887_call_ack_0, ack => d_block_daemon_CP_6409_elements(36)); -- 
    -- CP-element group 37:  join  fork  transition  input  output  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	29 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (14) 
      -- CP-element group 37: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12887_update_completed_
      -- CP-element group 37: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12887_Update/$exit
      -- CP-element group 37: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12887_Update/cca
      -- CP-element group 37: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12892_sample_start_
      -- CP-element group 37: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/R_K4_12888_sample_start_
      -- CP-element group 37: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/R_K4_12888_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/R_K4_12888_update_start_
      -- CP-element group 37: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/R_K4_12888_update_completed_
      -- CP-element group 37: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/R_RConstant_5_12889_sample_start_
      -- CP-element group 37: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/R_RConstant_5_12889_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/R_RConstant_5_12889_update_start_
      -- CP-element group 37: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/R_RConstant_5_12889_update_completed_
      -- CP-element group 37: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12892_Sample/$entry
      -- CP-element group 37: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12892_Sample/crr
      -- 
    cca_6657_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_12887_call_ack_1, ack => d_block_daemon_CP_6409_elements(37)); -- 
    crr_6673_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_6673_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_6409_elements(37), ack => call_stmt_12892_call_req_0); -- 
    -- CP-element group 38:  transition  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12892_sample_completed_
      -- CP-element group 38: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12892_Sample/$exit
      -- CP-element group 38: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12892_Sample/cra
      -- 
    cra_6674_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_12892_call_ack_0, ack => d_block_daemon_CP_6409_elements(38)); -- 
    -- CP-element group 39:  join  fork  transition  input  output  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	29 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	40 
    -- CP-element group 39:  members (14) 
      -- CP-element group 39: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12892_update_completed_
      -- CP-element group 39: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12892_Update/$exit
      -- CP-element group 39: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12892_Update/cca
      -- CP-element group 39: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12897_sample_start_
      -- CP-element group 39: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/R_K5_12893_sample_start_
      -- CP-element group 39: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/R_K5_12893_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/R_K5_12893_update_start_
      -- CP-element group 39: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/R_K5_12893_update_completed_
      -- CP-element group 39: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/R_RConstant_6_12894_sample_start_
      -- CP-element group 39: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/R_RConstant_6_12894_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/R_RConstant_6_12894_update_start_
      -- CP-element group 39: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/R_RConstant_6_12894_update_completed_
      -- CP-element group 39: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12897_Sample/$entry
      -- CP-element group 39: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12897_Sample/crr
      -- 
    cca_6679_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_12892_call_ack_1, ack => d_block_daemon_CP_6409_elements(39)); -- 
    crr_6695_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_6695_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_6409_elements(39), ack => call_stmt_12897_call_req_0); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	39 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12897_sample_completed_
      -- CP-element group 40: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12897_Sample/$exit
      -- CP-element group 40: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12897_Sample/cra
      -- 
    cra_6696_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_12897_call_ack_0, ack => d_block_daemon_CP_6409_elements(40)); -- 
    -- CP-element group 41:  join  fork  transition  input  output  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	29 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	42 
    -- CP-element group 41:  members (14) 
      -- CP-element group 41: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12897_update_completed_
      -- CP-element group 41: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12897_Update/$exit
      -- CP-element group 41: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12897_Update/cca
      -- CP-element group 41: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12902_sample_start_
      -- CP-element group 41: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/R_K6_12898_sample_start_
      -- CP-element group 41: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/R_K6_12898_sample_completed_
      -- CP-element group 41: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/R_K6_12898_update_start_
      -- CP-element group 41: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/R_K6_12898_update_completed_
      -- CP-element group 41: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/R_RConstant_7_12899_sample_start_
      -- CP-element group 41: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/R_RConstant_7_12899_sample_completed_
      -- CP-element group 41: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/R_RConstant_7_12899_update_start_
      -- CP-element group 41: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/R_RConstant_7_12899_update_completed_
      -- CP-element group 41: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12902_Sample/$entry
      -- CP-element group 41: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12902_Sample/crr
      -- 
    cca_6701_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_12897_call_ack_1, ack => d_block_daemon_CP_6409_elements(41)); -- 
    crr_6717_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_6717_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_6409_elements(41), ack => call_stmt_12902_call_req_0); -- 
    -- CP-element group 42:  transition  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	41 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12902_sample_completed_
      -- CP-element group 42: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12902_Sample/$exit
      -- CP-element group 42: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12902_Sample/cra
      -- 
    cra_6718_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_12902_call_ack_0, ack => d_block_daemon_CP_6409_elements(42)); -- 
    -- CP-element group 43:  join  fork  transition  input  output  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	29 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	44 
    -- CP-element group 43:  members (14) 
      -- CP-element group 43: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/R_RConstant_8_12904_update_start_
      -- CP-element group 43: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/R_K7_12903_update_completed_
      -- CP-element group 43: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12907_Sample/$entry
      -- CP-element group 43: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12907_Sample/crr
      -- CP-element group 43: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/R_RConstant_8_12904_update_completed_
      -- CP-element group 43: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/R_RConstant_8_12904_sample_start_
      -- CP-element group 43: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/R_RConstant_8_12904_sample_completed_
      -- CP-element group 43: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/R_K7_12903_update_start_
      -- CP-element group 43: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/R_K7_12903_sample_completed_
      -- CP-element group 43: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/R_K7_12903_sample_start_
      -- CP-element group 43: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12902_update_completed_
      -- CP-element group 43: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12902_Update/$exit
      -- CP-element group 43: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12902_Update/cca
      -- CP-element group 43: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12907_sample_start_
      -- 
    cca_6723_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_12902_call_ack_1, ack => d_block_daemon_CP_6409_elements(43)); -- 
    crr_6739_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_6739_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_6409_elements(43), ack => call_stmt_12907_call_req_0); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	43 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12907_Sample/cra
      -- CP-element group 44: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12907_Sample/$exit
      -- CP-element group 44: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12907_sample_completed_
      -- 
    cra_6740_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_12907_call_ack_0, ack => d_block_daemon_CP_6409_elements(44)); -- 
    -- CP-element group 45:  join  fork  transition  input  output  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	29 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45:  members (14) 
      -- CP-element group 45: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12907_Update/cca
      -- CP-element group 45: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12907_Update/$exit
      -- CP-element group 45: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12912_sample_start_
      -- CP-element group 45: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12907_update_completed_
      -- CP-element group 45: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12912_Sample/crr
      -- CP-element group 45: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12912_Sample/$entry
      -- CP-element group 45: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/R_RConstant_9_12909_update_completed_
      -- CP-element group 45: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/R_RConstant_9_12909_update_start_
      -- CP-element group 45: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/R_RConstant_9_12909_sample_completed_
      -- CP-element group 45: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/R_RConstant_9_12909_sample_start_
      -- CP-element group 45: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/R_K8_12908_update_completed_
      -- CP-element group 45: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/R_K8_12908_update_start_
      -- CP-element group 45: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/R_K8_12908_sample_completed_
      -- CP-element group 45: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/R_K8_12908_sample_start_
      -- 
    cca_6745_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_12907_call_ack_1, ack => d_block_daemon_CP_6409_elements(45)); -- 
    crr_6761_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_6761_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_6409_elements(45), ack => call_stmt_12912_call_req_0); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12912_Sample/cra
      -- CP-element group 46: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12912_Sample/$exit
      -- CP-element group 46: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12912_sample_completed_
      -- 
    cra_6762_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_12912_call_ack_0, ack => d_block_daemon_CP_6409_elements(46)); -- 
    -- CP-element group 47:  join  fork  transition  input  output  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	29 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	48 
    -- CP-element group 47:  members (14) 
      -- CP-element group 47: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/R_RConstant_10_12914_update_start_
      -- CP-element group 47: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/R_RConstant_10_12914_update_completed_
      -- CP-element group 47: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12917_Sample/$entry
      -- CP-element group 47: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12917_Sample/crr
      -- CP-element group 47: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12912_update_completed_
      -- CP-element group 47: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/R_RConstant_10_12914_sample_completed_
      -- CP-element group 47: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/R_RConstant_10_12914_sample_start_
      -- CP-element group 47: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/R_K9_12913_update_completed_
      -- CP-element group 47: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/R_K9_12913_update_start_
      -- CP-element group 47: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/R_K9_12913_sample_completed_
      -- CP-element group 47: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/R_K9_12913_sample_start_
      -- CP-element group 47: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12917_sample_start_
      -- CP-element group 47: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12912_Update/cca
      -- CP-element group 47: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12912_Update/$exit
      -- 
    cca_6767_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_12912_call_ack_1, ack => d_block_daemon_CP_6409_elements(47)); -- 
    crr_6783_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_6783_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_6409_elements(47), ack => call_stmt_12917_call_req_0); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	47 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12917_Sample/$exit
      -- CP-element group 48: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12917_Sample/cra
      -- CP-element group 48: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12917_sample_completed_
      -- 
    cra_6784_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_12917_call_ack_0, ack => d_block_daemon_CP_6409_elements(48)); -- 
    -- CP-element group 49:  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	29 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	8 
    -- CP-element group 49:  members (4) 
      -- CP-element group 49: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12917_Update/cca
      -- CP-element group 49: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12917_Update/$exit
      -- CP-element group 49: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/call_stmt_12917_update_completed_
      -- CP-element group 49: 	 branch_block_stmt_12832/call_stmt_12872_to_call_stmt_12917/$exit
      -- 
    cca_6789_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_12917_call_ack_1, ack => d_block_daemon_CP_6409_elements(49)); -- 
    -- CP-element group 50:  transition  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	9 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50:  members (1) 
      -- CP-element group 50: 	 branch_block_stmt_12832/do_while_stmt_12924/$entry
      -- 
    d_block_daemon_CP_6409_elements(50) <= d_block_daemon_CP_6409_elements(9);
    -- CP-element group 51:  place  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	57 
    -- CP-element group 51:  members (1) 
      -- CP-element group 51: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924__entry__
      -- 
    d_block_daemon_CP_6409_elements(51) <= d_block_daemon_CP_6409_elements(50);
    -- CP-element group 52:  merge  place  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	193 
    -- CP-element group 52:  members (1) 
      -- CP-element group 52: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924__exit__
      -- 
    -- Element group d_block_daemon_CP_6409_elements(52) is bound as output of CP function.
    -- CP-element group 53:  merge  place  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	56 
    -- CP-element group 53:  members (1) 
      -- CP-element group 53: 	 branch_block_stmt_12832/do_while_stmt_12924/loop_back
      -- 
    -- Element group d_block_daemon_CP_6409_elements(53) is bound as output of CP function.
    -- CP-element group 54:  branch  place  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	59 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	189 
    -- CP-element group 54: 	191 
    -- CP-element group 54:  members (1) 
      -- CP-element group 54: 	 branch_block_stmt_12832/do_while_stmt_12924/condition_done
      -- 
    d_block_daemon_CP_6409_elements(54) <= d_block_daemon_CP_6409_elements(59);
    -- CP-element group 55:  branch  place  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	249 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (1) 
      -- CP-element group 55: 	 branch_block_stmt_12832/do_while_stmt_12924/loop_body_done
      -- 
    d_block_daemon_CP_6409_elements(55) <= d_block_daemon_CP_6409_elements(249);
    -- CP-element group 56:  transition  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	53 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	64 
    -- CP-element group 56:  members (1) 
      -- CP-element group 56: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/back_edge_to_loop_body
      -- 
    d_block_daemon_CP_6409_elements(56) <= d_block_daemon_CP_6409_elements(53);
    -- CP-element group 57:  transition  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	51 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	66 
    -- CP-element group 57:  members (1) 
      -- CP-element group 57: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/first_time_through_loop_body
      -- 
    d_block_daemon_CP_6409_elements(57) <= d_block_daemon_CP_6409_elements(51);
    -- CP-element group 58:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	126 
    -- CP-element group 58: 	128 
    -- CP-element group 58: 	132 
    -- CP-element group 58: 	135 
    -- CP-element group 58: 	137 
    -- CP-element group 58: 	141 
    -- CP-element group 58: 	144 
    -- CP-element group 58: 	146 
    -- CP-element group 58: 	159 
    -- CP-element group 58: 	162 
    -- CP-element group 58: 	164 
    -- CP-element group 58: 	168 
    -- CP-element group 58: 	171 
    -- CP-element group 58: 	173 
    -- CP-element group 58: 	177 
    -- CP-element group 58: 	188 
    -- CP-element group 58: 	108 
    -- CP-element group 58: 	110 
    -- CP-element group 58: 	99 
    -- CP-element group 58: 	101 
    -- CP-element group 58: 	84 
    -- CP-element group 58: 	86 
    -- CP-element group 58: 	80 
    -- CP-element group 58: 	60 
    -- CP-element group 58: 	61 
    -- CP-element group 58: 	153 
    -- CP-element group 58: 	155 
    -- CP-element group 58: 	150 
    -- CP-element group 58: 	123 
    -- CP-element group 58: 	117 
    -- CP-element group 58: 	119 
    -- CP-element group 58: 	105 
    -- CP-element group 58: 	96 
    -- CP-element group 58: 	90 
    -- CP-element group 58: 	92 
    -- CP-element group 58: 	114 
    -- CP-element group 58:  members (28) 
      -- CP-element group 58: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_K9_12943_sample_completed_
      -- CP-element group 58: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_K9_12943_sample_start_
      -- CP-element group 58: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/loop_body_start
      -- CP-element group 58: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/$entry
      -- CP-element group 58: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_K10_12935_sample_completed_
      -- CP-element group 58: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_K10_12935_sample_start_
      -- CP-element group 58: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_K8_12951_sample_start_
      -- CP-element group 58: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_K8_12951_sample_completed_
      -- CP-element group 58: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_K7_12959_sample_start_
      -- CP-element group 58: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_K7_12959_sample_completed_
      -- CP-element group 58: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_K6_12967_sample_start_
      -- CP-element group 58: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_K6_12967_sample_completed_
      -- CP-element group 58: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_K5_12975_sample_start_
      -- CP-element group 58: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_K5_12975_sample_completed_
      -- CP-element group 58: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_K4_12983_sample_start_
      -- CP-element group 58: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_K4_12983_sample_completed_
      -- CP-element group 58: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_K3_12991_sample_start_
      -- CP-element group 58: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_K3_12991_sample_completed_
      -- CP-element group 58: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_K2_12999_sample_start_
      -- CP-element group 58: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_K2_12999_sample_completed_
      -- CP-element group 58: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_K1_13007_sample_start_
      -- CP-element group 58: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_K1_13007_sample_completed_
      -- CP-element group 58: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_K0_13015_sample_start_
      -- CP-element group 58: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_K0_13015_sample_completed_
      -- CP-element group 58: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_countB_13032_sample_start_
      -- CP-element group 58: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_countB_13032_sample_completed_
      -- CP-element group 58: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_countB_13032_update_start_
      -- CP-element group 58: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_countB_13032_update_completed_
      -- 
    -- Element group d_block_daemon_CP_6409_elements(58) is bound as output of CP function.
    -- CP-element group 59:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	188 
    -- CP-element group 59: 	61 
    -- CP-element group 59: 	62 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	54 
    -- CP-element group 59:  members (1) 
      -- CP-element group 59: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/condition_evaluated
      -- 
    condition_evaluated_6804_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_6804_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_6409_elements(59), ack => do_while_stmt_12924_branch_req_0); -- 
    d_block_daemon_cp_element_group_59: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 2,1 => 2,2 => 2);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "d_block_daemon_cp_element_group_59"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= d_block_daemon_CP_6409_elements(188) & d_block_daemon_CP_6409_elements(61) & d_block_daemon_CP_6409_elements(62);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => d_block_daemon_CP_6409_elements(59), clk => clk, reset => reset); --
    end block;
    -- CP-element group 60:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	58 
    -- CP-element group 60: marked-predecessors 
    -- CP-element group 60: 	187 
    -- CP-element group 60: 	62 
    -- CP-element group 60: successors 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/aggregated_phi_sample_req
      -- CP-element group 60: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/phi_stmt_12926_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/phi_stmt_12926_sample_start__ps
      -- 
    d_block_daemon_cp_element_group_60: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 2,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 34) := "d_block_daemon_cp_element_group_60"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= d_block_daemon_CP_6409_elements(58) & d_block_daemon_CP_6409_elements(187) & d_block_daemon_CP_6409_elements(62);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => d_block_daemon_CP_6409_elements(60), clk => clk, reset => reset); --
    end block;
    -- CP-element group 61:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	58 
    -- CP-element group 61: marked-predecessors 
    -- CP-element group 61: 	186 
    -- CP-element group 61: 	63 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	59 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/phi_stmt_12926_update_start__ps
      -- CP-element group 61: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/phi_stmt_12926_update_start_
      -- CP-element group 61: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/aggregated_phi_update_req
      -- 
    d_block_daemon_cp_element_group_61: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 2,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "d_block_daemon_cp_element_group_61"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= d_block_daemon_CP_6409_elements(58) & d_block_daemon_CP_6409_elements(186) & d_block_daemon_CP_6409_elements(63);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => d_block_daemon_CP_6409_elements(61), clk => clk, reset => reset); --
    end block;
    -- CP-element group 62:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	185 
    -- CP-element group 62: 	59 
    -- CP-element group 62: marked-successors 
    -- CP-element group 62: 	60 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/phi_stmt_12926_sample_completed__ps
      -- CP-element group 62: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/phi_stmt_12926_sample_completed_
      -- CP-element group 62: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/aggregated_phi_sample_ack
      -- 
    -- Element group d_block_daemon_CP_6409_elements(62) is bound as output of CP function.
    -- CP-element group 63:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	184 
    -- CP-element group 63: marked-successors 
    -- CP-element group 63: 	61 
    -- CP-element group 63:  members (7) 
      -- CP-element group 63: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/phi_stmt_12926_update_completed__ps
      -- CP-element group 63: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/phi_stmt_12926_update_completed_
      -- CP-element group 63: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/aggregated_phi_update_ack
      -- CP-element group 63: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_count_var_13026_sample_start_
      -- CP-element group 63: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_count_var_13026_sample_completed_
      -- CP-element group 63: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_count_var_13026_update_start_
      -- CP-element group 63: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_count_var_13026_update_completed_
      -- 
    -- Element group d_block_daemon_CP_6409_elements(63) is bound as output of CP function.
    -- CP-element group 64:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	56 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (1) 
      -- CP-element group 64: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/phi_stmt_12926_loopback_trigger
      -- 
    d_block_daemon_CP_6409_elements(64) <= d_block_daemon_CP_6409_elements(56);
    -- CP-element group 65:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	70 
    -- CP-element group 65:  members (1) 
      -- CP-element group 65: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/phi_stmt_12926_loopback_sample_req
      -- 
    phi_stmt_12926_loopback_sample_req_6819_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_12926_loopback_sample_req_6819_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_6409_elements(65), ack => phi_stmt_12926_req_1); -- 
    -- Element group d_block_daemon_CP_6409_elements(65) is bound as output of CP function.
    -- CP-element group 66:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	57 
    -- CP-element group 66: successors 
    -- CP-element group 66:  members (1) 
      -- CP-element group 66: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/phi_stmt_12926_entry_trigger
      -- 
    d_block_daemon_CP_6409_elements(66) <= d_block_daemon_CP_6409_elements(57);
    -- CP-element group 67:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	69 
    -- CP-element group 67:  members (1) 
      -- CP-element group 67: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/phi_stmt_12926_entry_sample_req
      -- 
    phi_stmt_12926_entry_sample_req_6821_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_12926_entry_sample_req_6821_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_6409_elements(67), ack => phi_stmt_12926_req_0); -- 
    -- Element group d_block_daemon_CP_6409_elements(67) is bound as output of CP function.
    -- CP-element group 68:  transition  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: successors 
    -- CP-element group 68:  members (1) 
      -- CP-element group 68: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/phi_stmt_12926_merged_reqs
      -- 
    -- Element group d_block_daemon_CP_6409_elements(68) is bound as output of CP function.
    -- CP-element group 69:  transition  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	67 
    -- CP-element group 69: successors 
    -- CP-element group 69:  members (1) 
      -- CP-element group 69: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/phi_stmt_12926_entry_sample_req__merge_in
      -- 
    d_block_daemon_CP_6409_elements(69) <= d_block_daemon_CP_6409_elements(67);
    -- CP-element group 70:  transition  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	65 
    -- CP-element group 70: successors 
    -- CP-element group 70:  members (1) 
      -- CP-element group 70: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/phi_stmt_12926_loopback_sample_req__merge_in
      -- 
    d_block_daemon_CP_6409_elements(70) <= d_block_daemon_CP_6409_elements(65);
    -- CP-element group 71:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	249 
    -- CP-element group 71:  members (1) 
      -- CP-element group 71: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/phi_stmt_12926_phi_mux_ack
      -- 
    phi_stmt_12926_phi_mux_ack_6826_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_12926_ack_0, ack => d_block_daemon_CP_6409_elements(71)); -- 
    -- CP-element group 72:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: successors 
    -- CP-element group 72:  members (4) 
      -- CP-element group 72: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_ZERO_COUNT_12928_sample_start_
      -- CP-element group 72: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_ZERO_COUNT_12928_sample_completed__ps
      -- CP-element group 72: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_ZERO_COUNT_12928_sample_start__ps
      -- CP-element group 72: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_ZERO_COUNT_12928_sample_completed_
      -- 
    -- Element group d_block_daemon_CP_6409_elements(72) is bound as output of CP function.
    -- CP-element group 73:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	75 
    -- CP-element group 73:  members (2) 
      -- CP-element group 73: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_ZERO_COUNT_12928_update_start__ps
      -- CP-element group 73: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_ZERO_COUNT_12928_update_start_
      -- 
    -- Element group d_block_daemon_CP_6409_elements(73) is bound as output of CP function.
    -- CP-element group 74:  join  transition  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	75 
    -- CP-element group 74: successors 
    -- CP-element group 74:  members (1) 
      -- CP-element group 74: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_ZERO_COUNT_12928_update_completed__ps
      -- 
    d_block_daemon_CP_6409_elements(74) <= d_block_daemon_CP_6409_elements(75);
    -- CP-element group 75:  transition  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	73 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	74 
    -- CP-element group 75:  members (1) 
      -- CP-element group 75: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_ZERO_COUNT_12928_update_completed_
      -- 
    -- Element group d_block_daemon_CP_6409_elements(75) is a control-delay.
    cp_element_75_delay: control_delay_element  generic map(name => " 75_delay", delay_value => 1)  port map(req => d_block_daemon_CP_6409_elements(73), ack => d_block_daemon_CP_6409_elements(75), clk => clk, reset =>reset);
    -- CP-element group 76:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	78 
    -- CP-element group 76:  members (4) 
      -- CP-element group 76: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_n_count_var_12929_Sample/req
      -- CP-element group 76: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_n_count_var_12929_Sample/$entry
      -- CP-element group 76: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_n_count_var_12929_sample_start_
      -- CP-element group 76: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_n_count_var_12929_sample_start__ps
      -- 
    req_6847_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6847_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_6409_elements(76), ack => n_count_var_13029_12929_buf_req_0); -- 
    -- Element group d_block_daemon_CP_6409_elements(76) is bound as output of CP function.
    -- CP-element group 77:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	79 
    -- CP-element group 77:  members (4) 
      -- CP-element group 77: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_n_count_var_12929_Update/req
      -- CP-element group 77: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_n_count_var_12929_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_n_count_var_12929_update_start_
      -- CP-element group 77: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_n_count_var_12929_update_start__ps
      -- 
    req_6852_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6852_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_6409_elements(77), ack => n_count_var_13029_12929_buf_req_1); -- 
    -- Element group d_block_daemon_CP_6409_elements(77) is bound as output of CP function.
    -- CP-element group 78:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	76 
    -- CP-element group 78: successors 
    -- CP-element group 78:  members (4) 
      -- CP-element group 78: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_n_count_var_12929_Sample/ack
      -- CP-element group 78: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_n_count_var_12929_Sample/$exit
      -- CP-element group 78: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_n_count_var_12929_sample_completed_
      -- CP-element group 78: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_n_count_var_12929_sample_completed__ps
      -- 
    ack_6848_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_count_var_13029_12929_buf_ack_0, ack => d_block_daemon_CP_6409_elements(78)); -- 
    -- CP-element group 79:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	77 
    -- CP-element group 79: successors 
    -- CP-element group 79:  members (4) 
      -- CP-element group 79: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_n_count_var_12929_Update/ack
      -- CP-element group 79: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_n_count_var_12929_Update/$exit
      -- CP-element group 79: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_n_count_var_12929_update_completed_
      -- CP-element group 79: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_n_count_var_12929_update_completed__ps
      -- 
    ack_6853_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_count_var_13029_12929_buf_ack_1, ack => d_block_daemon_CP_6409_elements(79)); -- 
    -- CP-element group 80:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	58 
    -- CP-element group 80: marked-predecessors 
    -- CP-element group 80: 	82 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	82 
    -- CP-element group 80:  members (3) 
      -- CP-element group 80: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/RPIPE_d_in_buf_12932_Sample/rr
      -- CP-element group 80: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/RPIPE_d_in_buf_12932_Sample/$entry
      -- CP-element group 80: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/RPIPE_d_in_buf_12932_sample_start_
      -- 
    rr_6862_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6862_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_6409_elements(80), ack => RPIPE_d_in_buf_12932_inst_req_0); -- 
    d_block_daemon_cp_element_group_80: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 2,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 34) := "d_block_daemon_cp_element_group_80"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= d_block_daemon_CP_6409_elements(58) & d_block_daemon_CP_6409_elements(82);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => d_block_daemon_CP_6409_elements(80), clk => clk, reset => reset); --
    end block;
    -- CP-element group 81:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	82 
    -- CP-element group 81: marked-predecessors 
    -- CP-element group 81: 	83 
    -- CP-element group 81: 	97 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	83 
    -- CP-element group 81:  members (3) 
      -- CP-element group 81: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/RPIPE_d_in_buf_12932_Update/$entry
      -- CP-element group 81: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/RPIPE_d_in_buf_12932_update_start_
      -- CP-element group 81: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/RPIPE_d_in_buf_12932_Update/cr
      -- 
    cr_6867_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6867_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_6409_elements(81), ack => RPIPE_d_in_buf_12932_inst_req_1); -- 
    d_block_daemon_cp_element_group_81: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 2,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "d_block_daemon_cp_element_group_81"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= d_block_daemon_CP_6409_elements(82) & d_block_daemon_CP_6409_elements(83) & d_block_daemon_CP_6409_elements(97);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => d_block_daemon_CP_6409_elements(81), clk => clk, reset => reset); --
    end block;
    -- CP-element group 82:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	80 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	81 
    -- CP-element group 82: marked-successors 
    -- CP-element group 82: 	80 
    -- CP-element group 82:  members (3) 
      -- CP-element group 82: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/RPIPE_d_in_buf_12932_Sample/ra
      -- CP-element group 82: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/RPIPE_d_in_buf_12932_Sample/$exit
      -- CP-element group 82: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/RPIPE_d_in_buf_12932_sample_completed_
      -- 
    ra_6863_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_d_in_buf_12932_inst_ack_0, ack => d_block_daemon_CP_6409_elements(82)); -- 
    -- CP-element group 83:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	81 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	89 
    -- CP-element group 83: marked-successors 
    -- CP-element group 83: 	81 
    -- CP-element group 83:  members (7) 
      -- CP-element group 83: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/RPIPE_d_in_buf_12932_update_completed_
      -- CP-element group 83: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_in128_12938_sample_completed_
      -- CP-element group 83: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_in128_12938_sample_start_
      -- CP-element group 83: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/RPIPE_d_in_buf_12932_Update/ca
      -- CP-element group 83: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_in128_12938_update_start_
      -- CP-element group 83: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/RPIPE_d_in_buf_12932_Update/$exit
      -- CP-element group 83: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_in128_12938_update_completed_
      -- 
    ca_6868_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_d_in_buf_12932_inst_ack_1, ack => d_block_daemon_CP_6409_elements(83)); -- 
    -- CP-element group 84:  join  transition  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	58 
    -- CP-element group 84: marked-predecessors 
    -- CP-element group 84: 	87 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	85 
    -- CP-element group 84:  members (2) 
      -- CP-element group 84: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_K10_12935_update_start_
      -- CP-element group 84: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_K10_12935_update_completed_
      -- 
    d_block_daemon_cp_element_group_84: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 2,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 34) := "d_block_daemon_cp_element_group_84"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= d_block_daemon_CP_6409_elements(58) & d_block_daemon_CP_6409_elements(87);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => d_block_daemon_CP_6409_elements(84), clk => clk, reset => reset); --
    end block;
    -- CP-element group 85:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	84 
    -- CP-element group 85: marked-predecessors 
    -- CP-element group 85: 	87 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	87 
    -- CP-element group 85:  members (3) 
      -- CP-element group 85: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_12936_Sample/req
      -- CP-element group 85: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_12936_Sample/$entry
      -- CP-element group 85: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_12936_sample_start_
      -- 
    req_6880_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6880_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_6409_elements(85), ack => W_K10_12936_delayed_1_12934_inst_req_0); -- 
    d_block_daemon_cp_element_group_85: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 2,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 34) := "d_block_daemon_cp_element_group_85"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= d_block_daemon_CP_6409_elements(84) & d_block_daemon_CP_6409_elements(87);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => d_block_daemon_CP_6409_elements(85), clk => clk, reset => reset); --
    end block;
    -- CP-element group 86:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	58 
    -- CP-element group 86: marked-predecessors 
    -- CP-element group 86: 	88 
    -- CP-element group 86: 	97 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	88 
    -- CP-element group 86:  members (3) 
      -- CP-element group 86: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_12936_Update/req
      -- CP-element group 86: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_12936_Update/$entry
      -- CP-element group 86: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_12936_update_start_
      -- 
    req_6885_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6885_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_6409_elements(86), ack => W_K10_12936_delayed_1_12934_inst_req_1); -- 
    d_block_daemon_cp_element_group_86: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 2,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "d_block_daemon_cp_element_group_86"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= d_block_daemon_CP_6409_elements(58) & d_block_daemon_CP_6409_elements(88) & d_block_daemon_CP_6409_elements(97);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => d_block_daemon_CP_6409_elements(86), clk => clk, reset => reset); --
    end block;
    -- CP-element group 87:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	85 
    -- CP-element group 87: successors 
    -- CP-element group 87: marked-successors 
    -- CP-element group 87: 	84 
    -- CP-element group 87: 	85 
    -- CP-element group 87:  members (3) 
      -- CP-element group 87: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_12936_Sample/ack
      -- CP-element group 87: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_12936_Sample/$exit
      -- CP-element group 87: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_12936_sample_completed_
      -- 
    ack_6881_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_K10_12936_delayed_1_12934_inst_ack_0, ack => d_block_daemon_CP_6409_elements(87)); -- 
    -- CP-element group 88:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	86 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	89 
    -- CP-element group 88: marked-successors 
    -- CP-element group 88: 	86 
    -- CP-element group 88:  members (7) 
      -- CP-element group 88: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_12936_Update/ack
      -- CP-element group 88: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_12936_Update/$exit
      -- CP-element group 88: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_K10_12936_delayed_1_12939_update_completed_
      -- CP-element group 88: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_K10_12936_delayed_1_12939_update_start_
      -- CP-element group 88: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_12936_update_completed_
      -- CP-element group 88: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_K10_12936_delayed_1_12939_sample_completed_
      -- CP-element group 88: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_K10_12936_delayed_1_12939_sample_start_
      -- 
    ack_6886_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_K10_12936_delayed_1_12934_inst_ack_1, ack => d_block_daemon_CP_6409_elements(88)); -- 
    -- CP-element group 89:  join  transition  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	83 
    -- CP-element group 89: 	88 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	95 
    -- CP-element group 89:  members (16) 
      -- CP-element group 89: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/XOR_u128_u128_12940_sample_completed_
      -- CP-element group 89: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/XOR_u128_u128_12940_Update/ca
      -- CP-element group 89: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/XOR_u128_u128_12940_sample_start_
      -- CP-element group 89: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/XOR_u128_u128_12940_Update/cr
      -- CP-element group 89: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/XOR_u128_u128_12940_Update/$exit
      -- CP-element group 89: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/XOR_u128_u128_12940_Update/$entry
      -- CP-element group 89: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/XOR_u128_u128_12940_Sample/ra
      -- CP-element group 89: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/XOR_u128_u128_12940_Sample/rr
      -- CP-element group 89: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/XOR_u128_u128_12940_Sample/$exit
      -- CP-element group 89: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/XOR_u128_u128_12940_Sample/$entry
      -- CP-element group 89: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_round_S10_12945_update_start_
      -- CP-element group 89: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_round_S10_12945_update_completed_
      -- CP-element group 89: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/XOR_u128_u128_12940_update_completed_
      -- CP-element group 89: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_round_S10_12945_sample_start_
      -- CP-element group 89: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_round_S10_12945_sample_completed_
      -- CP-element group 89: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/XOR_u128_u128_12940_update_start_
      -- 
    d_block_daemon_cp_element_group_89: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 2,1 => 2);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "d_block_daemon_cp_element_group_89"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= d_block_daemon_CP_6409_elements(83) & d_block_daemon_CP_6409_elements(88);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => d_block_daemon_CP_6409_elements(89), clk => clk, reset => reset); --
    end block;
    -- CP-element group 90:  join  transition  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	58 
    -- CP-element group 90: marked-predecessors 
    -- CP-element group 90: 	93 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	91 
    -- CP-element group 90:  members (2) 
      -- CP-element group 90: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_K9_12943_update_completed_
      -- CP-element group 90: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_K9_12943_update_start_
      -- 
    d_block_daemon_cp_element_group_90: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 2,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 34) := "d_block_daemon_cp_element_group_90"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= d_block_daemon_CP_6409_elements(58) & d_block_daemon_CP_6409_elements(93);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => d_block_daemon_CP_6409_elements(90), clk => clk, reset => reset); --
    end block;
    -- CP-element group 91:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	90 
    -- CP-element group 91: marked-predecessors 
    -- CP-element group 91: 	93 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	93 
    -- CP-element group 91:  members (3) 
      -- CP-element group 91: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_12944_Sample/req
      -- CP-element group 91: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_12944_sample_start_
      -- CP-element group 91: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_12944_Sample/$entry
      -- 
    req_6920_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6920_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_6409_elements(91), ack => W_K9_12940_delayed_1_12942_inst_req_0); -- 
    d_block_daemon_cp_element_group_91: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 2,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 34) := "d_block_daemon_cp_element_group_91"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= d_block_daemon_CP_6409_elements(90) & d_block_daemon_CP_6409_elements(93);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => d_block_daemon_CP_6409_elements(91), clk => clk, reset => reset); --
    end block;
    -- CP-element group 92:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	58 
    -- CP-element group 92: marked-predecessors 
    -- CP-element group 92: 	97 
    -- CP-element group 92: 	94 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	94 
    -- CP-element group 92:  members (3) 
      -- CP-element group 92: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_12944_Update/$entry
      -- CP-element group 92: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_12944_update_start_
      -- CP-element group 92: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_12944_Update/req
      -- 
    req_6925_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6925_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_6409_elements(92), ack => W_K9_12940_delayed_1_12942_inst_req_1); -- 
    d_block_daemon_cp_element_group_92: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 2,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "d_block_daemon_cp_element_group_92"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= d_block_daemon_CP_6409_elements(58) & d_block_daemon_CP_6409_elements(97) & d_block_daemon_CP_6409_elements(94);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => d_block_daemon_CP_6409_elements(92), clk => clk, reset => reset); --
    end block;
    -- CP-element group 93:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	91 
    -- CP-element group 93: successors 
    -- CP-element group 93: marked-successors 
    -- CP-element group 93: 	90 
    -- CP-element group 93: 	91 
    -- CP-element group 93:  members (3) 
      -- CP-element group 93: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_12944_Sample/$exit
      -- CP-element group 93: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_12944_Sample/ack
      -- CP-element group 93: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_12944_sample_completed_
      -- 
    ack_6921_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_K9_12940_delayed_1_12942_inst_ack_0, ack => d_block_daemon_CP_6409_elements(93)); -- 
    -- CP-element group 94:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	92 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	95 
    -- CP-element group 94: marked-successors 
    -- CP-element group 94: 	92 
    -- CP-element group 94:  members (7) 
      -- CP-element group 94: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_12944_update_completed_
      -- CP-element group 94: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_12944_Update/$exit
      -- CP-element group 94: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_12944_Update/ack
      -- CP-element group 94: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_K9_12940_delayed_1_12946_update_start_
      -- CP-element group 94: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_K9_12940_delayed_1_12946_update_completed_
      -- CP-element group 94: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_K9_12940_delayed_1_12946_sample_start_
      -- CP-element group 94: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_K9_12940_delayed_1_12946_sample_completed_
      -- 
    ack_6926_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_K9_12940_delayed_1_12942_inst_ack_1, ack => d_block_daemon_CP_6409_elements(94)); -- 
    -- CP-element group 95:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	89 
    -- CP-element group 95: 	94 
    -- CP-element group 95: marked-predecessors 
    -- CP-element group 95: 	97 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	97 
    -- CP-element group 95:  members (3) 
      -- CP-element group 95: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_12949_sample_start_
      -- CP-element group 95: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_12949_Sample/$entry
      -- CP-element group 95: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_12949_Sample/crr
      -- 
    crr_6942_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_6942_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_6409_elements(95), ack => call_stmt_12949_call_req_0); -- 
    d_block_daemon_cp_element_group_95: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 2,1 => 2,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 34) := "d_block_daemon_cp_element_group_95"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= d_block_daemon_CP_6409_elements(89) & d_block_daemon_CP_6409_elements(94) & d_block_daemon_CP_6409_elements(97);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => d_block_daemon_CP_6409_elements(95), clk => clk, reset => reset); --
    end block;
    -- CP-element group 96:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	58 
    -- CP-element group 96: marked-predecessors 
    -- CP-element group 96: 	106 
    -- CP-element group 96: 	98 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	98 
    -- CP-element group 96:  members (3) 
      -- CP-element group 96: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_12949_update_start_
      -- CP-element group 96: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_12949_Update/$entry
      -- CP-element group 96: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_12949_Update/ccr
      -- 
    ccr_6947_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_6947_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_6409_elements(96), ack => call_stmt_12949_call_req_1); -- 
    d_block_daemon_cp_element_group_96: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 2,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "d_block_daemon_cp_element_group_96"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= d_block_daemon_CP_6409_elements(58) & d_block_daemon_CP_6409_elements(106) & d_block_daemon_CP_6409_elements(98);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => d_block_daemon_CP_6409_elements(96), clk => clk, reset => reset); --
    end block;
    -- CP-element group 97:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	95 
    -- CP-element group 97: successors 
    -- CP-element group 97: marked-successors 
    -- CP-element group 97: 	86 
    -- CP-element group 97: 	81 
    -- CP-element group 97: 	95 
    -- CP-element group 97: 	92 
    -- CP-element group 97:  members (3) 
      -- CP-element group 97: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_12949_sample_completed_
      -- CP-element group 97: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_12949_Sample/$exit
      -- CP-element group 97: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_12949_Sample/cra
      -- 
    cra_6943_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_12949_call_ack_0, ack => d_block_daemon_CP_6409_elements(97)); -- 
    -- CP-element group 98:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	96 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	104 
    -- CP-element group 98: marked-successors 
    -- CP-element group 98: 	96 
    -- CP-element group 98:  members (7) 
      -- CP-element group 98: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_12949_update_completed_
      -- CP-element group 98: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_12949_Update/$exit
      -- CP-element group 98: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_12949_Update/cca
      -- CP-element group 98: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_round_S9_12953_sample_start_
      -- CP-element group 98: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_round_S9_12953_sample_completed_
      -- CP-element group 98: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_round_S9_12953_update_start_
      -- CP-element group 98: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_round_S9_12953_update_completed_
      -- 
    cca_6948_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_12949_call_ack_1, ack => d_block_daemon_CP_6409_elements(98)); -- 
    -- CP-element group 99:  join  transition  bypass  pipeline-parent 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	58 
    -- CP-element group 99: marked-predecessors 
    -- CP-element group 99: 	102 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	100 
    -- CP-element group 99:  members (2) 
      -- CP-element group 99: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_K8_12951_update_start_
      -- CP-element group 99: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_K8_12951_update_completed_
      -- 
    d_block_daemon_cp_element_group_99: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 2,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 34) := "d_block_daemon_cp_element_group_99"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= d_block_daemon_CP_6409_elements(58) & d_block_daemon_CP_6409_elements(102);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => d_block_daemon_CP_6409_elements(99), clk => clk, reset => reset); --
    end block;
    -- CP-element group 100:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	99 
    -- CP-element group 100: marked-predecessors 
    -- CP-element group 100: 	102 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	102 
    -- CP-element group 100:  members (3) 
      -- CP-element group 100: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_12952_sample_start_
      -- CP-element group 100: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_12952_Sample/$entry
      -- CP-element group 100: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_12952_Sample/req
      -- 
    req_6960_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6960_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_6409_elements(100), ack => W_K8_12945_delayed_2_12950_inst_req_0); -- 
    d_block_daemon_cp_element_group_100: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 2,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "d_block_daemon_cp_element_group_100"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= d_block_daemon_CP_6409_elements(99) & d_block_daemon_CP_6409_elements(102);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => d_block_daemon_CP_6409_elements(100), clk => clk, reset => reset); --
    end block;
    -- CP-element group 101:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	58 
    -- CP-element group 101: marked-predecessors 
    -- CP-element group 101: 	106 
    -- CP-element group 101: 	103 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	103 
    -- CP-element group 101:  members (3) 
      -- CP-element group 101: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_12952_update_start_
      -- CP-element group 101: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_12952_Update/$entry
      -- CP-element group 101: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_12952_Update/req
      -- 
    req_6965_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6965_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_6409_elements(101), ack => W_K8_12945_delayed_2_12950_inst_req_1); -- 
    d_block_daemon_cp_element_group_101: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 2,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "d_block_daemon_cp_element_group_101"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= d_block_daemon_CP_6409_elements(58) & d_block_daemon_CP_6409_elements(106) & d_block_daemon_CP_6409_elements(103);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => d_block_daemon_CP_6409_elements(101), clk => clk, reset => reset); --
    end block;
    -- CP-element group 102:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	100 
    -- CP-element group 102: successors 
    -- CP-element group 102: marked-successors 
    -- CP-element group 102: 	99 
    -- CP-element group 102: 	100 
    -- CP-element group 102:  members (3) 
      -- CP-element group 102: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_12952_sample_completed_
      -- CP-element group 102: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_12952_Sample/$exit
      -- CP-element group 102: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_12952_Sample/ack
      -- 
    ack_6961_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_K8_12945_delayed_2_12950_inst_ack_0, ack => d_block_daemon_CP_6409_elements(102)); -- 
    -- CP-element group 103:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	101 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	104 
    -- CP-element group 103: marked-successors 
    -- CP-element group 103: 	101 
    -- CP-element group 103:  members (7) 
      -- CP-element group 103: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_12952_update_completed_
      -- CP-element group 103: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_12952_Update/$exit
      -- CP-element group 103: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_12952_Update/ack
      -- CP-element group 103: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_K8_12945_delayed_2_12954_sample_start_
      -- CP-element group 103: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_K8_12945_delayed_2_12954_sample_completed_
      -- CP-element group 103: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_K8_12945_delayed_2_12954_update_start_
      -- CP-element group 103: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_K8_12945_delayed_2_12954_update_completed_
      -- 
    ack_6966_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_K8_12945_delayed_2_12950_inst_ack_1, ack => d_block_daemon_CP_6409_elements(103)); -- 
    -- CP-element group 104:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	98 
    -- CP-element group 104: 	103 
    -- CP-element group 104: marked-predecessors 
    -- CP-element group 104: 	106 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	106 
    -- CP-element group 104:  members (3) 
      -- CP-element group 104: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_12957_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_12957_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_12957_Sample/crr
      -- 
    crr_6982_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_6982_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_6409_elements(104), ack => call_stmt_12957_call_req_0); -- 
    d_block_daemon_cp_element_group_104: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 2,1 => 2,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 35) := "d_block_daemon_cp_element_group_104"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= d_block_daemon_CP_6409_elements(98) & d_block_daemon_CP_6409_elements(103) & d_block_daemon_CP_6409_elements(106);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => d_block_daemon_CP_6409_elements(104), clk => clk, reset => reset); --
    end block;
    -- CP-element group 105:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	58 
    -- CP-element group 105: marked-predecessors 
    -- CP-element group 105: 	107 
    -- CP-element group 105: 	115 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	107 
    -- CP-element group 105:  members (3) 
      -- CP-element group 105: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_12957_update_start_
      -- CP-element group 105: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_12957_Update/$entry
      -- CP-element group 105: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_12957_Update/ccr
      -- 
    ccr_6987_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_6987_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_6409_elements(105), ack => call_stmt_12957_call_req_1); -- 
    d_block_daemon_cp_element_group_105: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 2,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "d_block_daemon_cp_element_group_105"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= d_block_daemon_CP_6409_elements(58) & d_block_daemon_CP_6409_elements(107) & d_block_daemon_CP_6409_elements(115);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => d_block_daemon_CP_6409_elements(105), clk => clk, reset => reset); --
    end block;
    -- CP-element group 106:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	104 
    -- CP-element group 106: successors 
    -- CP-element group 106: marked-successors 
    -- CP-element group 106: 	101 
    -- CP-element group 106: 	104 
    -- CP-element group 106: 	96 
    -- CP-element group 106:  members (3) 
      -- CP-element group 106: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_12957_sample_completed_
      -- CP-element group 106: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_12957_Sample/$exit
      -- CP-element group 106: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_12957_Sample/cra
      -- 
    cra_6983_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_12957_call_ack_0, ack => d_block_daemon_CP_6409_elements(106)); -- 
    -- CP-element group 107:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	105 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	113 
    -- CP-element group 107: marked-successors 
    -- CP-element group 107: 	105 
    -- CP-element group 107:  members (7) 
      -- CP-element group 107: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_12957_update_completed_
      -- CP-element group 107: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_12957_Update/$exit
      -- CP-element group 107: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_12957_Update/cca
      -- CP-element group 107: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_round_S8_12961_sample_start_
      -- CP-element group 107: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_round_S8_12961_sample_completed_
      -- CP-element group 107: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_round_S8_12961_update_start_
      -- CP-element group 107: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_round_S8_12961_update_completed_
      -- 
    cca_6988_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_12957_call_ack_1, ack => d_block_daemon_CP_6409_elements(107)); -- 
    -- CP-element group 108:  join  transition  bypass  pipeline-parent 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	58 
    -- CP-element group 108: marked-predecessors 
    -- CP-element group 108: 	111 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	109 
    -- CP-element group 108:  members (2) 
      -- CP-element group 108: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_K7_12959_update_start_
      -- CP-element group 108: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_K7_12959_update_completed_
      -- 
    d_block_daemon_cp_element_group_108: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 2,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "d_block_daemon_cp_element_group_108"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= d_block_daemon_CP_6409_elements(58) & d_block_daemon_CP_6409_elements(111);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => d_block_daemon_CP_6409_elements(108), clk => clk, reset => reset); --
    end block;
    -- CP-element group 109:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	108 
    -- CP-element group 109: marked-predecessors 
    -- CP-element group 109: 	111 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	111 
    -- CP-element group 109:  members (3) 
      -- CP-element group 109: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_12960_Sample/$entry
      -- CP-element group 109: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_12960_sample_start_
      -- CP-element group 109: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_12960_Sample/req
      -- 
    req_7000_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7000_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_6409_elements(109), ack => W_K7_12950_delayed_3_12958_inst_req_0); -- 
    d_block_daemon_cp_element_group_109: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 2,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "d_block_daemon_cp_element_group_109"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= d_block_daemon_CP_6409_elements(108) & d_block_daemon_CP_6409_elements(111);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => d_block_daemon_CP_6409_elements(109), clk => clk, reset => reset); --
    end block;
    -- CP-element group 110:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	58 
    -- CP-element group 110: marked-predecessors 
    -- CP-element group 110: 	115 
    -- CP-element group 110: 	112 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	112 
    -- CP-element group 110:  members (3) 
      -- CP-element group 110: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_12960_update_start_
      -- CP-element group 110: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_12960_Update/$entry
      -- CP-element group 110: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_12960_Update/req
      -- 
    req_7005_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7005_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_6409_elements(110), ack => W_K7_12950_delayed_3_12958_inst_req_1); -- 
    d_block_daemon_cp_element_group_110: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 2,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "d_block_daemon_cp_element_group_110"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= d_block_daemon_CP_6409_elements(58) & d_block_daemon_CP_6409_elements(115) & d_block_daemon_CP_6409_elements(112);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => d_block_daemon_CP_6409_elements(110), clk => clk, reset => reset); --
    end block;
    -- CP-element group 111:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	109 
    -- CP-element group 111: successors 
    -- CP-element group 111: marked-successors 
    -- CP-element group 111: 	108 
    -- CP-element group 111: 	109 
    -- CP-element group 111:  members (3) 
      -- CP-element group 111: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_12960_sample_completed_
      -- CP-element group 111: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_12960_Sample/$exit
      -- CP-element group 111: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_12960_Sample/ack
      -- 
    ack_7001_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_K7_12950_delayed_3_12958_inst_ack_0, ack => d_block_daemon_CP_6409_elements(111)); -- 
    -- CP-element group 112:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	110 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	113 
    -- CP-element group 112: marked-successors 
    -- CP-element group 112: 	110 
    -- CP-element group 112:  members (7) 
      -- CP-element group 112: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_12960_update_completed_
      -- CP-element group 112: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_12960_Update/$exit
      -- CP-element group 112: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_12960_Update/ack
      -- CP-element group 112: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_K7_12950_delayed_3_12962_sample_start_
      -- CP-element group 112: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_K7_12950_delayed_3_12962_sample_completed_
      -- CP-element group 112: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_K7_12950_delayed_3_12962_update_start_
      -- CP-element group 112: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_K7_12950_delayed_3_12962_update_completed_
      -- 
    ack_7006_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_K7_12950_delayed_3_12958_inst_ack_1, ack => d_block_daemon_CP_6409_elements(112)); -- 
    -- CP-element group 113:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	107 
    -- CP-element group 113: 	112 
    -- CP-element group 113: marked-predecessors 
    -- CP-element group 113: 	115 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	115 
    -- CP-element group 113:  members (3) 
      -- CP-element group 113: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_12965_sample_start_
      -- CP-element group 113: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_12965_Sample/$entry
      -- CP-element group 113: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_12965_Sample/crr
      -- 
    crr_7022_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_7022_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_6409_elements(113), ack => call_stmt_12965_call_req_0); -- 
    d_block_daemon_cp_element_group_113: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 2,1 => 2,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 35) := "d_block_daemon_cp_element_group_113"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= d_block_daemon_CP_6409_elements(107) & d_block_daemon_CP_6409_elements(112) & d_block_daemon_CP_6409_elements(115);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => d_block_daemon_CP_6409_elements(113), clk => clk, reset => reset); --
    end block;
    -- CP-element group 114:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	58 
    -- CP-element group 114: marked-predecessors 
    -- CP-element group 114: 	124 
    -- CP-element group 114: 	116 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	116 
    -- CP-element group 114:  members (3) 
      -- CP-element group 114: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_12965_update_start_
      -- CP-element group 114: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_12965_Update/$entry
      -- CP-element group 114: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_12965_Update/ccr
      -- 
    ccr_7027_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_7027_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_6409_elements(114), ack => call_stmt_12965_call_req_1); -- 
    d_block_daemon_cp_element_group_114: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 2,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "d_block_daemon_cp_element_group_114"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= d_block_daemon_CP_6409_elements(58) & d_block_daemon_CP_6409_elements(124) & d_block_daemon_CP_6409_elements(116);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => d_block_daemon_CP_6409_elements(114), clk => clk, reset => reset); --
    end block;
    -- CP-element group 115:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	113 
    -- CP-element group 115: successors 
    -- CP-element group 115: marked-successors 
    -- CP-element group 115: 	110 
    -- CP-element group 115: 	105 
    -- CP-element group 115: 	113 
    -- CP-element group 115:  members (3) 
      -- CP-element group 115: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_12965_sample_completed_
      -- CP-element group 115: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_12965_Sample/$exit
      -- CP-element group 115: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_12965_Sample/cra
      -- 
    cra_7023_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_12965_call_ack_0, ack => d_block_daemon_CP_6409_elements(115)); -- 
    -- CP-element group 116:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	114 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	122 
    -- CP-element group 116: marked-successors 
    -- CP-element group 116: 	114 
    -- CP-element group 116:  members (7) 
      -- CP-element group 116: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_12965_update_completed_
      -- CP-element group 116: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_12965_Update/$exit
      -- CP-element group 116: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_12965_Update/cca
      -- CP-element group 116: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_round_S7_12969_sample_start_
      -- CP-element group 116: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_round_S7_12969_sample_completed_
      -- CP-element group 116: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_round_S7_12969_update_start_
      -- CP-element group 116: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_round_S7_12969_update_completed_
      -- 
    cca_7028_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_12965_call_ack_1, ack => d_block_daemon_CP_6409_elements(116)); -- 
    -- CP-element group 117:  join  transition  bypass  pipeline-parent 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	58 
    -- CP-element group 117: marked-predecessors 
    -- CP-element group 117: 	120 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	118 
    -- CP-element group 117:  members (2) 
      -- CP-element group 117: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_K6_12967_update_start_
      -- CP-element group 117: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_K6_12967_update_completed_
      -- 
    d_block_daemon_cp_element_group_117: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 2,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "d_block_daemon_cp_element_group_117"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= d_block_daemon_CP_6409_elements(58) & d_block_daemon_CP_6409_elements(120);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => d_block_daemon_CP_6409_elements(117), clk => clk, reset => reset); --
    end block;
    -- CP-element group 118:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	117 
    -- CP-element group 118: marked-predecessors 
    -- CP-element group 118: 	120 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	120 
    -- CP-element group 118:  members (3) 
      -- CP-element group 118: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_12968_sample_start_
      -- CP-element group 118: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_12968_Sample/$entry
      -- CP-element group 118: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_12968_Sample/req
      -- 
    req_7040_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7040_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_6409_elements(118), ack => W_K6_12955_delayed_4_12966_inst_req_0); -- 
    d_block_daemon_cp_element_group_118: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 2,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "d_block_daemon_cp_element_group_118"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= d_block_daemon_CP_6409_elements(117) & d_block_daemon_CP_6409_elements(120);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => d_block_daemon_CP_6409_elements(118), clk => clk, reset => reset); --
    end block;
    -- CP-element group 119:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	58 
    -- CP-element group 119: marked-predecessors 
    -- CP-element group 119: 	124 
    -- CP-element group 119: 	121 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	121 
    -- CP-element group 119:  members (3) 
      -- CP-element group 119: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_12968_update_start_
      -- CP-element group 119: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_12968_Update/$entry
      -- CP-element group 119: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_12968_Update/req
      -- 
    req_7045_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7045_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_6409_elements(119), ack => W_K6_12955_delayed_4_12966_inst_req_1); -- 
    d_block_daemon_cp_element_group_119: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 2,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "d_block_daemon_cp_element_group_119"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= d_block_daemon_CP_6409_elements(58) & d_block_daemon_CP_6409_elements(124) & d_block_daemon_CP_6409_elements(121);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => d_block_daemon_CP_6409_elements(119), clk => clk, reset => reset); --
    end block;
    -- CP-element group 120:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	118 
    -- CP-element group 120: successors 
    -- CP-element group 120: marked-successors 
    -- CP-element group 120: 	117 
    -- CP-element group 120: 	118 
    -- CP-element group 120:  members (3) 
      -- CP-element group 120: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_12968_sample_completed_
      -- CP-element group 120: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_12968_Sample/$exit
      -- CP-element group 120: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_12968_Sample/ack
      -- 
    ack_7041_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_K6_12955_delayed_4_12966_inst_ack_0, ack => d_block_daemon_CP_6409_elements(120)); -- 
    -- CP-element group 121:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	119 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	122 
    -- CP-element group 121: marked-successors 
    -- CP-element group 121: 	119 
    -- CP-element group 121:  members (7) 
      -- CP-element group 121: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_12968_update_completed_
      -- CP-element group 121: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_12968_Update/$exit
      -- CP-element group 121: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_12968_Update/ack
      -- CP-element group 121: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_K6_12955_delayed_4_12970_sample_start_
      -- CP-element group 121: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_K6_12955_delayed_4_12970_sample_completed_
      -- CP-element group 121: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_K6_12955_delayed_4_12970_update_start_
      -- CP-element group 121: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_K6_12955_delayed_4_12970_update_completed_
      -- 
    ack_7046_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_K6_12955_delayed_4_12966_inst_ack_1, ack => d_block_daemon_CP_6409_elements(121)); -- 
    -- CP-element group 122:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	121 
    -- CP-element group 122: 	116 
    -- CP-element group 122: marked-predecessors 
    -- CP-element group 122: 	124 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	124 
    -- CP-element group 122:  members (3) 
      -- CP-element group 122: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_12973_sample_start_
      -- CP-element group 122: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_12973_Sample/$entry
      -- CP-element group 122: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_12973_Sample/crr
      -- 
    crr_7062_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_7062_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_6409_elements(122), ack => call_stmt_12973_call_req_0); -- 
    d_block_daemon_cp_element_group_122: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 2,1 => 2,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 35) := "d_block_daemon_cp_element_group_122"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= d_block_daemon_CP_6409_elements(121) & d_block_daemon_CP_6409_elements(116) & d_block_daemon_CP_6409_elements(124);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => d_block_daemon_CP_6409_elements(122), clk => clk, reset => reset); --
    end block;
    -- CP-element group 123:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	58 
    -- CP-element group 123: marked-predecessors 
    -- CP-element group 123: 	125 
    -- CP-element group 123: 	133 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	125 
    -- CP-element group 123:  members (3) 
      -- CP-element group 123: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_12973_update_start_
      -- CP-element group 123: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_12973_Update/$entry
      -- CP-element group 123: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_12973_Update/ccr
      -- 
    ccr_7067_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_7067_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_6409_elements(123), ack => call_stmt_12973_call_req_1); -- 
    d_block_daemon_cp_element_group_123: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 2,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "d_block_daemon_cp_element_group_123"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= d_block_daemon_CP_6409_elements(58) & d_block_daemon_CP_6409_elements(125) & d_block_daemon_CP_6409_elements(133);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => d_block_daemon_CP_6409_elements(123), clk => clk, reset => reset); --
    end block;
    -- CP-element group 124:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	122 
    -- CP-element group 124: successors 
    -- CP-element group 124: marked-successors 
    -- CP-element group 124: 	122 
    -- CP-element group 124: 	119 
    -- CP-element group 124: 	114 
    -- CP-element group 124:  members (3) 
      -- CP-element group 124: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_12973_sample_completed_
      -- CP-element group 124: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_12973_Sample/$exit
      -- CP-element group 124: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_12973_Sample/cra
      -- 
    cra_7063_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_12973_call_ack_0, ack => d_block_daemon_CP_6409_elements(124)); -- 
    -- CP-element group 125:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	123 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	131 
    -- CP-element group 125: marked-successors 
    -- CP-element group 125: 	123 
    -- CP-element group 125:  members (7) 
      -- CP-element group 125: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_12973_update_completed_
      -- CP-element group 125: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_12973_Update/$exit
      -- CP-element group 125: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_12973_Update/cca
      -- CP-element group 125: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_round_S6_12977_sample_start_
      -- CP-element group 125: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_round_S6_12977_sample_completed_
      -- CP-element group 125: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_round_S6_12977_update_start_
      -- CP-element group 125: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_round_S6_12977_update_completed_
      -- 
    cca_7068_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_12973_call_ack_1, ack => d_block_daemon_CP_6409_elements(125)); -- 
    -- CP-element group 126:  join  transition  bypass  pipeline-parent 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	58 
    -- CP-element group 126: marked-predecessors 
    -- CP-element group 126: 	129 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	127 
    -- CP-element group 126:  members (2) 
      -- CP-element group 126: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_K5_12975_update_start_
      -- CP-element group 126: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_K5_12975_update_completed_
      -- 
    d_block_daemon_cp_element_group_126: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 2,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "d_block_daemon_cp_element_group_126"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= d_block_daemon_CP_6409_elements(58) & d_block_daemon_CP_6409_elements(129);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => d_block_daemon_CP_6409_elements(126), clk => clk, reset => reset); --
    end block;
    -- CP-element group 127:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	126 
    -- CP-element group 127: marked-predecessors 
    -- CP-element group 127: 	129 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	129 
    -- CP-element group 127:  members (3) 
      -- CP-element group 127: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_12976_sample_start_
      -- CP-element group 127: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_12976_Sample/$entry
      -- CP-element group 127: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_12976_Sample/req
      -- 
    req_7080_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7080_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_6409_elements(127), ack => W_K5_12960_delayed_5_12974_inst_req_0); -- 
    d_block_daemon_cp_element_group_127: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 2,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "d_block_daemon_cp_element_group_127"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= d_block_daemon_CP_6409_elements(126) & d_block_daemon_CP_6409_elements(129);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => d_block_daemon_CP_6409_elements(127), clk => clk, reset => reset); --
    end block;
    -- CP-element group 128:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	58 
    -- CP-element group 128: marked-predecessors 
    -- CP-element group 128: 	130 
    -- CP-element group 128: 	133 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	130 
    -- CP-element group 128:  members (3) 
      -- CP-element group 128: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_12976_update_start_
      -- CP-element group 128: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_12976_Update/$entry
      -- CP-element group 128: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_12976_Update/req
      -- 
    req_7085_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7085_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_6409_elements(128), ack => W_K5_12960_delayed_5_12974_inst_req_1); -- 
    d_block_daemon_cp_element_group_128: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 2,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "d_block_daemon_cp_element_group_128"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= d_block_daemon_CP_6409_elements(58) & d_block_daemon_CP_6409_elements(130) & d_block_daemon_CP_6409_elements(133);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => d_block_daemon_CP_6409_elements(128), clk => clk, reset => reset); --
    end block;
    -- CP-element group 129:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	127 
    -- CP-element group 129: successors 
    -- CP-element group 129: marked-successors 
    -- CP-element group 129: 	126 
    -- CP-element group 129: 	127 
    -- CP-element group 129:  members (3) 
      -- CP-element group 129: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_12976_sample_completed_
      -- CP-element group 129: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_12976_Sample/$exit
      -- CP-element group 129: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_12976_Sample/ack
      -- 
    ack_7081_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 129_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_K5_12960_delayed_5_12974_inst_ack_0, ack => d_block_daemon_CP_6409_elements(129)); -- 
    -- CP-element group 130:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	128 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	131 
    -- CP-element group 130: marked-successors 
    -- CP-element group 130: 	128 
    -- CP-element group 130:  members (7) 
      -- CP-element group 130: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_12976_update_completed_
      -- CP-element group 130: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_12976_Update/$exit
      -- CP-element group 130: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_12976_Update/ack
      -- CP-element group 130: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_K5_12960_delayed_5_12978_sample_start_
      -- CP-element group 130: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_K5_12960_delayed_5_12978_sample_completed_
      -- CP-element group 130: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_K5_12960_delayed_5_12978_update_start_
      -- CP-element group 130: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_K5_12960_delayed_5_12978_update_completed_
      -- 
    ack_7086_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 130_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_K5_12960_delayed_5_12974_inst_ack_1, ack => d_block_daemon_CP_6409_elements(130)); -- 
    -- CP-element group 131:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	125 
    -- CP-element group 131: 	130 
    -- CP-element group 131: marked-predecessors 
    -- CP-element group 131: 	133 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	133 
    -- CP-element group 131:  members (3) 
      -- CP-element group 131: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_12981_sample_start_
      -- CP-element group 131: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_12981_Sample/$entry
      -- CP-element group 131: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_12981_Sample/crr
      -- 
    crr_7102_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_7102_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_6409_elements(131), ack => call_stmt_12981_call_req_0); -- 
    d_block_daemon_cp_element_group_131: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 2,1 => 2,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 35) := "d_block_daemon_cp_element_group_131"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= d_block_daemon_CP_6409_elements(125) & d_block_daemon_CP_6409_elements(130) & d_block_daemon_CP_6409_elements(133);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => d_block_daemon_CP_6409_elements(131), clk => clk, reset => reset); --
    end block;
    -- CP-element group 132:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	58 
    -- CP-element group 132: marked-predecessors 
    -- CP-element group 132: 	134 
    -- CP-element group 132: 	142 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	134 
    -- CP-element group 132:  members (3) 
      -- CP-element group 132: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_12981_update_start_
      -- CP-element group 132: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_12981_Update/$entry
      -- CP-element group 132: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_12981_Update/ccr
      -- 
    ccr_7107_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_7107_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_6409_elements(132), ack => call_stmt_12981_call_req_1); -- 
    d_block_daemon_cp_element_group_132: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 2,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "d_block_daemon_cp_element_group_132"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= d_block_daemon_CP_6409_elements(58) & d_block_daemon_CP_6409_elements(134) & d_block_daemon_CP_6409_elements(142);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => d_block_daemon_CP_6409_elements(132), clk => clk, reset => reset); --
    end block;
    -- CP-element group 133:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	131 
    -- CP-element group 133: successors 
    -- CP-element group 133: marked-successors 
    -- CP-element group 133: 	128 
    -- CP-element group 133: 	131 
    -- CP-element group 133: 	123 
    -- CP-element group 133:  members (3) 
      -- CP-element group 133: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_12981_sample_completed_
      -- CP-element group 133: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_12981_Sample/$exit
      -- CP-element group 133: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_12981_Sample/cra
      -- 
    cra_7103_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_12981_call_ack_0, ack => d_block_daemon_CP_6409_elements(133)); -- 
    -- CP-element group 134:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	132 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	140 
    -- CP-element group 134: marked-successors 
    -- CP-element group 134: 	132 
    -- CP-element group 134:  members (7) 
      -- CP-element group 134: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_12981_update_completed_
      -- CP-element group 134: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_12981_Update/$exit
      -- CP-element group 134: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_12981_Update/cca
      -- CP-element group 134: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_round_S5_12985_sample_start_
      -- CP-element group 134: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_round_S5_12985_sample_completed_
      -- CP-element group 134: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_round_S5_12985_update_start_
      -- CP-element group 134: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_round_S5_12985_update_completed_
      -- 
    cca_7108_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 134_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_12981_call_ack_1, ack => d_block_daemon_CP_6409_elements(134)); -- 
    -- CP-element group 135:  join  transition  bypass  pipeline-parent 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	58 
    -- CP-element group 135: marked-predecessors 
    -- CP-element group 135: 	138 
    -- CP-element group 135: successors 
    -- CP-element group 135: 	136 
    -- CP-element group 135:  members (2) 
      -- CP-element group 135: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_K4_12983_update_start_
      -- CP-element group 135: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_K4_12983_update_completed_
      -- 
    d_block_daemon_cp_element_group_135: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 2,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "d_block_daemon_cp_element_group_135"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= d_block_daemon_CP_6409_elements(58) & d_block_daemon_CP_6409_elements(138);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => d_block_daemon_CP_6409_elements(135), clk => clk, reset => reset); --
    end block;
    -- CP-element group 136:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	135 
    -- CP-element group 136: marked-predecessors 
    -- CP-element group 136: 	138 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	138 
    -- CP-element group 136:  members (3) 
      -- CP-element group 136: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_12984_sample_start_
      -- CP-element group 136: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_12984_Sample/$entry
      -- CP-element group 136: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_12984_Sample/req
      -- 
    req_7120_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7120_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_6409_elements(136), ack => W_K4_12965_delayed_6_12982_inst_req_0); -- 
    d_block_daemon_cp_element_group_136: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 2,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "d_block_daemon_cp_element_group_136"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= d_block_daemon_CP_6409_elements(135) & d_block_daemon_CP_6409_elements(138);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => d_block_daemon_CP_6409_elements(136), clk => clk, reset => reset); --
    end block;
    -- CP-element group 137:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	58 
    -- CP-element group 137: marked-predecessors 
    -- CP-element group 137: 	139 
    -- CP-element group 137: 	142 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	139 
    -- CP-element group 137:  members (3) 
      -- CP-element group 137: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_12984_update_start_
      -- CP-element group 137: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_12984_Update/$entry
      -- CP-element group 137: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_12984_Update/req
      -- 
    req_7125_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7125_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_6409_elements(137), ack => W_K4_12965_delayed_6_12982_inst_req_1); -- 
    d_block_daemon_cp_element_group_137: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 2,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "d_block_daemon_cp_element_group_137"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= d_block_daemon_CP_6409_elements(58) & d_block_daemon_CP_6409_elements(139) & d_block_daemon_CP_6409_elements(142);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => d_block_daemon_CP_6409_elements(137), clk => clk, reset => reset); --
    end block;
    -- CP-element group 138:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	136 
    -- CP-element group 138: successors 
    -- CP-element group 138: marked-successors 
    -- CP-element group 138: 	135 
    -- CP-element group 138: 	136 
    -- CP-element group 138:  members (3) 
      -- CP-element group 138: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_12984_sample_completed_
      -- CP-element group 138: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_12984_Sample/$exit
      -- CP-element group 138: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_12984_Sample/ack
      -- 
    ack_7121_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 138_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_K4_12965_delayed_6_12982_inst_ack_0, ack => d_block_daemon_CP_6409_elements(138)); -- 
    -- CP-element group 139:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	137 
    -- CP-element group 139: successors 
    -- CP-element group 139: 	140 
    -- CP-element group 139: marked-successors 
    -- CP-element group 139: 	137 
    -- CP-element group 139:  members (7) 
      -- CP-element group 139: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_12984_update_completed_
      -- CP-element group 139: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_12984_Update/$exit
      -- CP-element group 139: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_12984_Update/ack
      -- CP-element group 139: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_K4_12965_delayed_6_12986_sample_start_
      -- CP-element group 139: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_K4_12965_delayed_6_12986_sample_completed_
      -- CP-element group 139: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_K4_12965_delayed_6_12986_update_start_
      -- CP-element group 139: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_K4_12965_delayed_6_12986_update_completed_
      -- 
    ack_7126_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 139_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_K4_12965_delayed_6_12982_inst_ack_1, ack => d_block_daemon_CP_6409_elements(139)); -- 
    -- CP-element group 140:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	134 
    -- CP-element group 140: 	139 
    -- CP-element group 140: marked-predecessors 
    -- CP-element group 140: 	142 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	142 
    -- CP-element group 140:  members (3) 
      -- CP-element group 140: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_12989_sample_start_
      -- CP-element group 140: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_12989_Sample/$entry
      -- CP-element group 140: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_12989_Sample/crr
      -- 
    crr_7142_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_7142_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_6409_elements(140), ack => call_stmt_12989_call_req_0); -- 
    d_block_daemon_cp_element_group_140: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 2,1 => 2,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 35) := "d_block_daemon_cp_element_group_140"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= d_block_daemon_CP_6409_elements(134) & d_block_daemon_CP_6409_elements(139) & d_block_daemon_CP_6409_elements(142);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => d_block_daemon_CP_6409_elements(140), clk => clk, reset => reset); --
    end block;
    -- CP-element group 141:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	58 
    -- CP-element group 141: marked-predecessors 
    -- CP-element group 141: 	143 
    -- CP-element group 141: 	151 
    -- CP-element group 141: successors 
    -- CP-element group 141: 	143 
    -- CP-element group 141:  members (3) 
      -- CP-element group 141: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_12989_update_start_
      -- CP-element group 141: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_12989_Update/$entry
      -- CP-element group 141: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_12989_Update/ccr
      -- 
    ccr_7147_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_7147_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_6409_elements(141), ack => call_stmt_12989_call_req_1); -- 
    d_block_daemon_cp_element_group_141: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 2,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "d_block_daemon_cp_element_group_141"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= d_block_daemon_CP_6409_elements(58) & d_block_daemon_CP_6409_elements(143) & d_block_daemon_CP_6409_elements(151);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => d_block_daemon_CP_6409_elements(141), clk => clk, reset => reset); --
    end block;
    -- CP-element group 142:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	140 
    -- CP-element group 142: successors 
    -- CP-element group 142: marked-successors 
    -- CP-element group 142: 	132 
    -- CP-element group 142: 	137 
    -- CP-element group 142: 	140 
    -- CP-element group 142:  members (3) 
      -- CP-element group 142: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_12989_sample_completed_
      -- CP-element group 142: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_12989_Sample/$exit
      -- CP-element group 142: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_12989_Sample/cra
      -- 
    cra_7143_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 142_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_12989_call_ack_0, ack => d_block_daemon_CP_6409_elements(142)); -- 
    -- CP-element group 143:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	141 
    -- CP-element group 143: successors 
    -- CP-element group 143: 	149 
    -- CP-element group 143: marked-successors 
    -- CP-element group 143: 	141 
    -- CP-element group 143:  members (7) 
      -- CP-element group 143: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_12989_update_completed_
      -- CP-element group 143: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_12989_Update/$exit
      -- CP-element group 143: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_12989_Update/cca
      -- CP-element group 143: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_round_S4_12993_sample_start_
      -- CP-element group 143: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_round_S4_12993_sample_completed_
      -- CP-element group 143: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_round_S4_12993_update_start_
      -- CP-element group 143: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_round_S4_12993_update_completed_
      -- 
    cca_7148_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 143_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_12989_call_ack_1, ack => d_block_daemon_CP_6409_elements(143)); -- 
    -- CP-element group 144:  join  transition  bypass  pipeline-parent 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	58 
    -- CP-element group 144: marked-predecessors 
    -- CP-element group 144: 	147 
    -- CP-element group 144: successors 
    -- CP-element group 144: 	145 
    -- CP-element group 144:  members (2) 
      -- CP-element group 144: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_K3_12991_update_start_
      -- CP-element group 144: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_K3_12991_update_completed_
      -- 
    d_block_daemon_cp_element_group_144: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 2,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "d_block_daemon_cp_element_group_144"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= d_block_daemon_CP_6409_elements(58) & d_block_daemon_CP_6409_elements(147);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => d_block_daemon_CP_6409_elements(144), clk => clk, reset => reset); --
    end block;
    -- CP-element group 145:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	144 
    -- CP-element group 145: marked-predecessors 
    -- CP-element group 145: 	147 
    -- CP-element group 145: successors 
    -- CP-element group 145: 	147 
    -- CP-element group 145:  members (3) 
      -- CP-element group 145: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_12992_sample_start_
      -- CP-element group 145: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_12992_Sample/$entry
      -- CP-element group 145: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_12992_Sample/req
      -- 
    req_7160_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7160_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_6409_elements(145), ack => W_K3_12970_delayed_7_12990_inst_req_0); -- 
    d_block_daemon_cp_element_group_145: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 2,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "d_block_daemon_cp_element_group_145"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= d_block_daemon_CP_6409_elements(144) & d_block_daemon_CP_6409_elements(147);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => d_block_daemon_CP_6409_elements(145), clk => clk, reset => reset); --
    end block;
    -- CP-element group 146:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	58 
    -- CP-element group 146: marked-predecessors 
    -- CP-element group 146: 	151 
    -- CP-element group 146: 	148 
    -- CP-element group 146: successors 
    -- CP-element group 146: 	148 
    -- CP-element group 146:  members (3) 
      -- CP-element group 146: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_12992_update_start_
      -- CP-element group 146: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_12992_Update/$entry
      -- CP-element group 146: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_12992_Update/req
      -- 
    req_7165_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7165_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_6409_elements(146), ack => W_K3_12970_delayed_7_12990_inst_req_1); -- 
    d_block_daemon_cp_element_group_146: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 2,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "d_block_daemon_cp_element_group_146"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= d_block_daemon_CP_6409_elements(58) & d_block_daemon_CP_6409_elements(151) & d_block_daemon_CP_6409_elements(148);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => d_block_daemon_CP_6409_elements(146), clk => clk, reset => reset); --
    end block;
    -- CP-element group 147:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	145 
    -- CP-element group 147: successors 
    -- CP-element group 147: marked-successors 
    -- CP-element group 147: 	144 
    -- CP-element group 147: 	145 
    -- CP-element group 147:  members (3) 
      -- CP-element group 147: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_12992_sample_completed_
      -- CP-element group 147: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_12992_Sample/$exit
      -- CP-element group 147: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_12992_Sample/ack
      -- 
    ack_7161_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 147_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_K3_12970_delayed_7_12990_inst_ack_0, ack => d_block_daemon_CP_6409_elements(147)); -- 
    -- CP-element group 148:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	146 
    -- CP-element group 148: successors 
    -- CP-element group 148: 	149 
    -- CP-element group 148: marked-successors 
    -- CP-element group 148: 	146 
    -- CP-element group 148:  members (7) 
      -- CP-element group 148: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_12992_update_completed_
      -- CP-element group 148: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_12992_Update/$exit
      -- CP-element group 148: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_12992_Update/ack
      -- CP-element group 148: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_K3_12970_delayed_7_12994_sample_start_
      -- CP-element group 148: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_K3_12970_delayed_7_12994_sample_completed_
      -- CP-element group 148: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_K3_12970_delayed_7_12994_update_start_
      -- CP-element group 148: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_K3_12970_delayed_7_12994_update_completed_
      -- 
    ack_7166_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 148_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_K3_12970_delayed_7_12990_inst_ack_1, ack => d_block_daemon_CP_6409_elements(148)); -- 
    -- CP-element group 149:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	143 
    -- CP-element group 149: 	148 
    -- CP-element group 149: marked-predecessors 
    -- CP-element group 149: 	151 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	151 
    -- CP-element group 149:  members (3) 
      -- CP-element group 149: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_12997_sample_start_
      -- CP-element group 149: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_12997_Sample/$entry
      -- CP-element group 149: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_12997_Sample/crr
      -- 
    crr_7182_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_7182_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_6409_elements(149), ack => call_stmt_12997_call_req_0); -- 
    d_block_daemon_cp_element_group_149: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 2,1 => 2,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 35) := "d_block_daemon_cp_element_group_149"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= d_block_daemon_CP_6409_elements(143) & d_block_daemon_CP_6409_elements(148) & d_block_daemon_CP_6409_elements(151);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => d_block_daemon_CP_6409_elements(149), clk => clk, reset => reset); --
    end block;
    -- CP-element group 150:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	58 
    -- CP-element group 150: marked-predecessors 
    -- CP-element group 150: 	160 
    -- CP-element group 150: 	152 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	152 
    -- CP-element group 150:  members (3) 
      -- CP-element group 150: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_12997_update_start_
      -- CP-element group 150: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_12997_Update/$entry
      -- CP-element group 150: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_12997_Update/ccr
      -- 
    ccr_7187_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_7187_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_6409_elements(150), ack => call_stmt_12997_call_req_1); -- 
    d_block_daemon_cp_element_group_150: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 2,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "d_block_daemon_cp_element_group_150"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= d_block_daemon_CP_6409_elements(58) & d_block_daemon_CP_6409_elements(160) & d_block_daemon_CP_6409_elements(152);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => d_block_daemon_CP_6409_elements(150), clk => clk, reset => reset); --
    end block;
    -- CP-element group 151:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	149 
    -- CP-element group 151: successors 
    -- CP-element group 151: marked-successors 
    -- CP-element group 151: 	141 
    -- CP-element group 151: 	146 
    -- CP-element group 151: 	149 
    -- CP-element group 151:  members (3) 
      -- CP-element group 151: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_12997_sample_completed_
      -- CP-element group 151: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_12997_Sample/$exit
      -- CP-element group 151: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_12997_Sample/cra
      -- 
    cra_7183_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 151_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_12997_call_ack_0, ack => d_block_daemon_CP_6409_elements(151)); -- 
    -- CP-element group 152:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	150 
    -- CP-element group 152: successors 
    -- CP-element group 152: 	158 
    -- CP-element group 152: marked-successors 
    -- CP-element group 152: 	150 
    -- CP-element group 152:  members (7) 
      -- CP-element group 152: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_round_S3_13001_update_start_
      -- CP-element group 152: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_round_S3_13001_update_completed_
      -- CP-element group 152: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_12997_update_completed_
      -- CP-element group 152: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_12997_Update/$exit
      -- CP-element group 152: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_12997_Update/cca
      -- CP-element group 152: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_round_S3_13001_sample_start_
      -- CP-element group 152: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_round_S3_13001_sample_completed_
      -- 
    cca_7188_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_12997_call_ack_1, ack => d_block_daemon_CP_6409_elements(152)); -- 
    -- CP-element group 153:  join  transition  bypass  pipeline-parent 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	58 
    -- CP-element group 153: marked-predecessors 
    -- CP-element group 153: 	156 
    -- CP-element group 153: successors 
    -- CP-element group 153: 	154 
    -- CP-element group 153:  members (2) 
      -- CP-element group 153: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_K2_12999_update_start_
      -- CP-element group 153: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_K2_12999_update_completed_
      -- 
    d_block_daemon_cp_element_group_153: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 2,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "d_block_daemon_cp_element_group_153"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= d_block_daemon_CP_6409_elements(58) & d_block_daemon_CP_6409_elements(156);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => d_block_daemon_CP_6409_elements(153), clk => clk, reset => reset); --
    end block;
    -- CP-element group 154:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	153 
    -- CP-element group 154: marked-predecessors 
    -- CP-element group 154: 	156 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	156 
    -- CP-element group 154:  members (3) 
      -- CP-element group 154: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_13000_sample_start_
      -- CP-element group 154: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_13000_Sample/$entry
      -- CP-element group 154: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_13000_Sample/req
      -- 
    req_7200_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7200_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_6409_elements(154), ack => W_K2_12975_delayed_8_12998_inst_req_0); -- 
    d_block_daemon_cp_element_group_154: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 2,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "d_block_daemon_cp_element_group_154"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= d_block_daemon_CP_6409_elements(153) & d_block_daemon_CP_6409_elements(156);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => d_block_daemon_CP_6409_elements(154), clk => clk, reset => reset); --
    end block;
    -- CP-element group 155:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	58 
    -- CP-element group 155: marked-predecessors 
    -- CP-element group 155: 	157 
    -- CP-element group 155: 	160 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	157 
    -- CP-element group 155:  members (3) 
      -- CP-element group 155: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_13000_update_start_
      -- CP-element group 155: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_13000_Update/$entry
      -- CP-element group 155: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_13000_Update/req
      -- 
    req_7205_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7205_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_6409_elements(155), ack => W_K2_12975_delayed_8_12998_inst_req_1); -- 
    d_block_daemon_cp_element_group_155: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 2,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "d_block_daemon_cp_element_group_155"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= d_block_daemon_CP_6409_elements(58) & d_block_daemon_CP_6409_elements(157) & d_block_daemon_CP_6409_elements(160);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => d_block_daemon_CP_6409_elements(155), clk => clk, reset => reset); --
    end block;
    -- CP-element group 156:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	154 
    -- CP-element group 156: successors 
    -- CP-element group 156: marked-successors 
    -- CP-element group 156: 	153 
    -- CP-element group 156: 	154 
    -- CP-element group 156:  members (3) 
      -- CP-element group 156: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_13000_sample_completed_
      -- CP-element group 156: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_13000_Sample/$exit
      -- CP-element group 156: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_13000_Sample/ack
      -- 
    ack_7201_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 156_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_K2_12975_delayed_8_12998_inst_ack_0, ack => d_block_daemon_CP_6409_elements(156)); -- 
    -- CP-element group 157:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	155 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	158 
    -- CP-element group 157: marked-successors 
    -- CP-element group 157: 	155 
    -- CP-element group 157:  members (7) 
      -- CP-element group 157: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_13000_update_completed_
      -- CP-element group 157: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_13000_Update/$exit
      -- CP-element group 157: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_13000_Update/ack
      -- CP-element group 157: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_K2_12975_delayed_8_13002_sample_start_
      -- CP-element group 157: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_K2_12975_delayed_8_13002_sample_completed_
      -- CP-element group 157: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_K2_12975_delayed_8_13002_update_start_
      -- CP-element group 157: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_K2_12975_delayed_8_13002_update_completed_
      -- 
    ack_7206_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 157_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_K2_12975_delayed_8_12998_inst_ack_1, ack => d_block_daemon_CP_6409_elements(157)); -- 
    -- CP-element group 158:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	157 
    -- CP-element group 158: 	152 
    -- CP-element group 158: marked-predecessors 
    -- CP-element group 158: 	160 
    -- CP-element group 158: successors 
    -- CP-element group 158: 	160 
    -- CP-element group 158:  members (3) 
      -- CP-element group 158: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_13005_sample_start_
      -- CP-element group 158: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_13005_Sample/$entry
      -- CP-element group 158: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_13005_Sample/crr
      -- 
    crr_7222_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_7222_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_6409_elements(158), ack => call_stmt_13005_call_req_0); -- 
    d_block_daemon_cp_element_group_158: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 2,1 => 2,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 35) := "d_block_daemon_cp_element_group_158"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= d_block_daemon_CP_6409_elements(157) & d_block_daemon_CP_6409_elements(152) & d_block_daemon_CP_6409_elements(160);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => d_block_daemon_CP_6409_elements(158), clk => clk, reset => reset); --
    end block;
    -- CP-element group 159:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	58 
    -- CP-element group 159: marked-predecessors 
    -- CP-element group 159: 	161 
    -- CP-element group 159: 	169 
    -- CP-element group 159: successors 
    -- CP-element group 159: 	161 
    -- CP-element group 159:  members (3) 
      -- CP-element group 159: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_13005_update_start_
      -- CP-element group 159: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_13005_Update/$entry
      -- CP-element group 159: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_13005_Update/ccr
      -- 
    ccr_7227_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_7227_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_6409_elements(159), ack => call_stmt_13005_call_req_1); -- 
    d_block_daemon_cp_element_group_159: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 2,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "d_block_daemon_cp_element_group_159"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= d_block_daemon_CP_6409_elements(58) & d_block_daemon_CP_6409_elements(161) & d_block_daemon_CP_6409_elements(169);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => d_block_daemon_CP_6409_elements(159), clk => clk, reset => reset); --
    end block;
    -- CP-element group 160:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	158 
    -- CP-element group 160: successors 
    -- CP-element group 160: marked-successors 
    -- CP-element group 160: 	158 
    -- CP-element group 160: 	155 
    -- CP-element group 160: 	150 
    -- CP-element group 160:  members (3) 
      -- CP-element group 160: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_13005_sample_completed_
      -- CP-element group 160: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_13005_Sample/$exit
      -- CP-element group 160: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_13005_Sample/cra
      -- 
    cra_7223_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 160_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_13005_call_ack_0, ack => d_block_daemon_CP_6409_elements(160)); -- 
    -- CP-element group 161:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	159 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	167 
    -- CP-element group 161: marked-successors 
    -- CP-element group 161: 	159 
    -- CP-element group 161:  members (7) 
      -- CP-element group 161: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_13005_update_completed_
      -- CP-element group 161: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_13005_Update/$exit
      -- CP-element group 161: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_13005_Update/cca
      -- CP-element group 161: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_round_S2_13009_sample_start_
      -- CP-element group 161: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_round_S2_13009_sample_completed_
      -- CP-element group 161: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_round_S2_13009_update_start_
      -- CP-element group 161: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_round_S2_13009_update_completed_
      -- 
    cca_7228_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 161_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_13005_call_ack_1, ack => d_block_daemon_CP_6409_elements(161)); -- 
    -- CP-element group 162:  join  transition  bypass  pipeline-parent 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	58 
    -- CP-element group 162: marked-predecessors 
    -- CP-element group 162: 	165 
    -- CP-element group 162: successors 
    -- CP-element group 162: 	163 
    -- CP-element group 162:  members (2) 
      -- CP-element group 162: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_K1_13007_update_start_
      -- CP-element group 162: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_K1_13007_update_completed_
      -- 
    d_block_daemon_cp_element_group_162: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 2,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "d_block_daemon_cp_element_group_162"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= d_block_daemon_CP_6409_elements(58) & d_block_daemon_CP_6409_elements(165);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => d_block_daemon_CP_6409_elements(162), clk => clk, reset => reset); --
    end block;
    -- CP-element group 163:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	162 
    -- CP-element group 163: marked-predecessors 
    -- CP-element group 163: 	165 
    -- CP-element group 163: successors 
    -- CP-element group 163: 	165 
    -- CP-element group 163:  members (3) 
      -- CP-element group 163: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_13008_sample_start_
      -- CP-element group 163: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_13008_Sample/$entry
      -- CP-element group 163: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_13008_Sample/req
      -- 
    req_7240_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7240_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_6409_elements(163), ack => W_K1_12980_delayed_9_13006_inst_req_0); -- 
    d_block_daemon_cp_element_group_163: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 2,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "d_block_daemon_cp_element_group_163"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= d_block_daemon_CP_6409_elements(162) & d_block_daemon_CP_6409_elements(165);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => d_block_daemon_CP_6409_elements(163), clk => clk, reset => reset); --
    end block;
    -- CP-element group 164:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: 	58 
    -- CP-element group 164: marked-predecessors 
    -- CP-element group 164: 	166 
    -- CP-element group 164: 	169 
    -- CP-element group 164: successors 
    -- CP-element group 164: 	166 
    -- CP-element group 164:  members (3) 
      -- CP-element group 164: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_13008_update_start_
      -- CP-element group 164: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_13008_Update/$entry
      -- CP-element group 164: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_13008_Update/req
      -- 
    req_7245_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7245_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_6409_elements(164), ack => W_K1_12980_delayed_9_13006_inst_req_1); -- 
    d_block_daemon_cp_element_group_164: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 2,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "d_block_daemon_cp_element_group_164"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= d_block_daemon_CP_6409_elements(58) & d_block_daemon_CP_6409_elements(166) & d_block_daemon_CP_6409_elements(169);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => d_block_daemon_CP_6409_elements(164), clk => clk, reset => reset); --
    end block;
    -- CP-element group 165:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	163 
    -- CP-element group 165: successors 
    -- CP-element group 165: marked-successors 
    -- CP-element group 165: 	162 
    -- CP-element group 165: 	163 
    -- CP-element group 165:  members (3) 
      -- CP-element group 165: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_13008_sample_completed_
      -- CP-element group 165: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_13008_Sample/$exit
      -- CP-element group 165: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_13008_Sample/ack
      -- 
    ack_7241_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 165_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_K1_12980_delayed_9_13006_inst_ack_0, ack => d_block_daemon_CP_6409_elements(165)); -- 
    -- CP-element group 166:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	164 
    -- CP-element group 166: successors 
    -- CP-element group 166: 	167 
    -- CP-element group 166: marked-successors 
    -- CP-element group 166: 	164 
    -- CP-element group 166:  members (7) 
      -- CP-element group 166: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_13008_update_completed_
      -- CP-element group 166: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_13008_Update/$exit
      -- CP-element group 166: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_13008_Update/ack
      -- CP-element group 166: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_K1_12980_delayed_9_13010_sample_start_
      -- CP-element group 166: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_K1_12980_delayed_9_13010_sample_completed_
      -- CP-element group 166: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_K1_12980_delayed_9_13010_update_start_
      -- CP-element group 166: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_K1_12980_delayed_9_13010_update_completed_
      -- 
    ack_7246_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 166_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_K1_12980_delayed_9_13006_inst_ack_1, ack => d_block_daemon_CP_6409_elements(166)); -- 
    -- CP-element group 167:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	161 
    -- CP-element group 167: 	166 
    -- CP-element group 167: marked-predecessors 
    -- CP-element group 167: 	169 
    -- CP-element group 167: successors 
    -- CP-element group 167: 	169 
    -- CP-element group 167:  members (3) 
      -- CP-element group 167: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_13013_sample_start_
      -- CP-element group 167: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_13013_Sample/$entry
      -- CP-element group 167: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_13013_Sample/crr
      -- 
    crr_7262_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_7262_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_6409_elements(167), ack => call_stmt_13013_call_req_0); -- 
    d_block_daemon_cp_element_group_167: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 2,1 => 2,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 35) := "d_block_daemon_cp_element_group_167"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= d_block_daemon_CP_6409_elements(161) & d_block_daemon_CP_6409_elements(166) & d_block_daemon_CP_6409_elements(169);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => d_block_daemon_CP_6409_elements(167), clk => clk, reset => reset); --
    end block;
    -- CP-element group 168:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	58 
    -- CP-element group 168: marked-predecessors 
    -- CP-element group 168: 	170 
    -- CP-element group 168: 	178 
    -- CP-element group 168: successors 
    -- CP-element group 168: 	170 
    -- CP-element group 168:  members (3) 
      -- CP-element group 168: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_13013_update_start_
      -- CP-element group 168: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_13013_Update/$entry
      -- CP-element group 168: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_13013_Update/ccr
      -- 
    ccr_7267_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_7267_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_6409_elements(168), ack => call_stmt_13013_call_req_1); -- 
    d_block_daemon_cp_element_group_168: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 2,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "d_block_daemon_cp_element_group_168"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= d_block_daemon_CP_6409_elements(58) & d_block_daemon_CP_6409_elements(170) & d_block_daemon_CP_6409_elements(178);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => d_block_daemon_CP_6409_elements(168), clk => clk, reset => reset); --
    end block;
    -- CP-element group 169:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	167 
    -- CP-element group 169: successors 
    -- CP-element group 169: marked-successors 
    -- CP-element group 169: 	159 
    -- CP-element group 169: 	164 
    -- CP-element group 169: 	167 
    -- CP-element group 169:  members (3) 
      -- CP-element group 169: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_13013_sample_completed_
      -- CP-element group 169: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_13013_Sample/$exit
      -- CP-element group 169: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_13013_Sample/cra
      -- 
    cra_7263_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 169_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_13013_call_ack_0, ack => d_block_daemon_CP_6409_elements(169)); -- 
    -- CP-element group 170:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	168 
    -- CP-element group 170: successors 
    -- CP-element group 170: 	176 
    -- CP-element group 170: marked-successors 
    -- CP-element group 170: 	168 
    -- CP-element group 170:  members (7) 
      -- CP-element group 170: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_13013_update_completed_
      -- CP-element group 170: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_13013_Update/$exit
      -- CP-element group 170: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_13013_Update/cca
      -- CP-element group 170: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_round_S1_13017_sample_start_
      -- CP-element group 170: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_round_S1_13017_sample_completed_
      -- CP-element group 170: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_round_S1_13017_update_start_
      -- CP-element group 170: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_round_S1_13017_update_completed_
      -- 
    cca_7268_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 170_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_13013_call_ack_1, ack => d_block_daemon_CP_6409_elements(170)); -- 
    -- CP-element group 171:  join  transition  bypass  pipeline-parent 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	58 
    -- CP-element group 171: marked-predecessors 
    -- CP-element group 171: 	174 
    -- CP-element group 171: successors 
    -- CP-element group 171: 	172 
    -- CP-element group 171:  members (2) 
      -- CP-element group 171: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_K0_13015_update_start_
      -- CP-element group 171: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_K0_13015_update_completed_
      -- 
    d_block_daemon_cp_element_group_171: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 2,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "d_block_daemon_cp_element_group_171"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= d_block_daemon_CP_6409_elements(58) & d_block_daemon_CP_6409_elements(174);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => d_block_daemon_CP_6409_elements(171), clk => clk, reset => reset); --
    end block;
    -- CP-element group 172:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	171 
    -- CP-element group 172: marked-predecessors 
    -- CP-element group 172: 	174 
    -- CP-element group 172: successors 
    -- CP-element group 172: 	174 
    -- CP-element group 172:  members (3) 
      -- CP-element group 172: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_13016_sample_start_
      -- CP-element group 172: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_13016_Sample/$entry
      -- CP-element group 172: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_13016_Sample/req
      -- 
    req_7280_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7280_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_6409_elements(172), ack => W_K0_12985_delayed_10_13014_inst_req_0); -- 
    d_block_daemon_cp_element_group_172: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 2,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "d_block_daemon_cp_element_group_172"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= d_block_daemon_CP_6409_elements(171) & d_block_daemon_CP_6409_elements(174);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => d_block_daemon_CP_6409_elements(172), clk => clk, reset => reset); --
    end block;
    -- CP-element group 173:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	58 
    -- CP-element group 173: marked-predecessors 
    -- CP-element group 173: 	175 
    -- CP-element group 173: 	178 
    -- CP-element group 173: successors 
    -- CP-element group 173: 	175 
    -- CP-element group 173:  members (3) 
      -- CP-element group 173: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_13016_update_start_
      -- CP-element group 173: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_13016_Update/$entry
      -- CP-element group 173: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_13016_Update/req
      -- 
    req_7285_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7285_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_6409_elements(173), ack => W_K0_12985_delayed_10_13014_inst_req_1); -- 
    d_block_daemon_cp_element_group_173: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 2,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "d_block_daemon_cp_element_group_173"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= d_block_daemon_CP_6409_elements(58) & d_block_daemon_CP_6409_elements(175) & d_block_daemon_CP_6409_elements(178);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => d_block_daemon_CP_6409_elements(173), clk => clk, reset => reset); --
    end block;
    -- CP-element group 174:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	172 
    -- CP-element group 174: successors 
    -- CP-element group 174: marked-successors 
    -- CP-element group 174: 	171 
    -- CP-element group 174: 	172 
    -- CP-element group 174:  members (3) 
      -- CP-element group 174: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_13016_sample_completed_
      -- CP-element group 174: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_13016_Sample/$exit
      -- CP-element group 174: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_13016_Sample/ack
      -- 
    ack_7281_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 174_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_K0_12985_delayed_10_13014_inst_ack_0, ack => d_block_daemon_CP_6409_elements(174)); -- 
    -- CP-element group 175:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	173 
    -- CP-element group 175: successors 
    -- CP-element group 175: 	176 
    -- CP-element group 175: marked-successors 
    -- CP-element group 175: 	173 
    -- CP-element group 175:  members (7) 
      -- CP-element group 175: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_13016_update_completed_
      -- CP-element group 175: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_13016_Update/$exit
      -- CP-element group 175: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/assign_stmt_13016_Update/ack
      -- CP-element group 175: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_K0_12985_delayed_10_13018_sample_start_
      -- CP-element group 175: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_K0_12985_delayed_10_13018_sample_completed_
      -- CP-element group 175: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_K0_12985_delayed_10_13018_update_start_
      -- CP-element group 175: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_K0_12985_delayed_10_13018_update_completed_
      -- 
    ack_7286_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 175_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_K0_12985_delayed_10_13014_inst_ack_1, ack => d_block_daemon_CP_6409_elements(175)); -- 
    -- CP-element group 176:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: 	170 
    -- CP-element group 176: 	175 
    -- CP-element group 176: marked-predecessors 
    -- CP-element group 176: 	178 
    -- CP-element group 176: successors 
    -- CP-element group 176: 	178 
    -- CP-element group 176:  members (3) 
      -- CP-element group 176: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_13021_sample_start_
      -- CP-element group 176: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_13021_Sample/$entry
      -- CP-element group 176: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_13021_Sample/crr
      -- 
    crr_7302_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_7302_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_6409_elements(176), ack => call_stmt_13021_call_req_0); -- 
    d_block_daemon_cp_element_group_176: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 2,1 => 2,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 35) := "d_block_daemon_cp_element_group_176"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= d_block_daemon_CP_6409_elements(170) & d_block_daemon_CP_6409_elements(175) & d_block_daemon_CP_6409_elements(178);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => d_block_daemon_CP_6409_elements(176), clk => clk, reset => reset); --
    end block;
    -- CP-element group 177:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	58 
    -- CP-element group 177: marked-predecessors 
    -- CP-element group 177: 	179 
    -- CP-element group 177: 	182 
    -- CP-element group 177: successors 
    -- CP-element group 177: 	179 
    -- CP-element group 177:  members (3) 
      -- CP-element group 177: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_13021_update_start_
      -- CP-element group 177: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_13021_Update/$entry
      -- CP-element group 177: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_13021_Update/ccr
      -- 
    ccr_7307_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_7307_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_6409_elements(177), ack => call_stmt_13021_call_req_1); -- 
    d_block_daemon_cp_element_group_177: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 2,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "d_block_daemon_cp_element_group_177"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= d_block_daemon_CP_6409_elements(58) & d_block_daemon_CP_6409_elements(179) & d_block_daemon_CP_6409_elements(182);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => d_block_daemon_CP_6409_elements(177), clk => clk, reset => reset); --
    end block;
    -- CP-element group 178:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	176 
    -- CP-element group 178: successors 
    -- CP-element group 178: marked-successors 
    -- CP-element group 178: 	168 
    -- CP-element group 178: 	173 
    -- CP-element group 178: 	176 
    -- CP-element group 178:  members (3) 
      -- CP-element group 178: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_13021_sample_completed_
      -- CP-element group 178: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_13021_Sample/$exit
      -- CP-element group 178: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_13021_Sample/cra
      -- 
    cra_7303_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 178_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_13021_call_ack_0, ack => d_block_daemon_CP_6409_elements(178)); -- 
    -- CP-element group 179:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	177 
    -- CP-element group 179: successors 
    -- CP-element group 179: 	180 
    -- CP-element group 179: marked-successors 
    -- CP-element group 179: 	177 
    -- CP-element group 179:  members (7) 
      -- CP-element group 179: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_13021_update_completed_
      -- CP-element group 179: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_13021_Update/$exit
      -- CP-element group 179: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/call_stmt_13021_Update/cca
      -- CP-element group 179: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_round_S0_13023_sample_start_
      -- CP-element group 179: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_round_S0_13023_sample_completed_
      -- CP-element group 179: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_round_S0_13023_update_start_
      -- CP-element group 179: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_round_S0_13023_update_completed_
      -- 
    cca_7308_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 179_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_13021_call_ack_1, ack => d_block_daemon_CP_6409_elements(179)); -- 
    -- CP-element group 180:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	179 
    -- CP-element group 180: marked-predecessors 
    -- CP-element group 180: 	182 
    -- CP-element group 180: successors 
    -- CP-element group 180: 	182 
    -- CP-element group 180:  members (3) 
      -- CP-element group 180: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/WPIPE_d_out_buf_13022_sample_start_
      -- CP-element group 180: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/WPIPE_d_out_buf_13022_Sample/$entry
      -- CP-element group 180: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/WPIPE_d_out_buf_13022_Sample/req
      -- 
    req_7320_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7320_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_6409_elements(180), ack => WPIPE_d_out_buf_13022_inst_req_0); -- 
    d_block_daemon_cp_element_group_180: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 2,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "d_block_daemon_cp_element_group_180"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= d_block_daemon_CP_6409_elements(179) & d_block_daemon_CP_6409_elements(182);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => d_block_daemon_CP_6409_elements(180), clk => clk, reset => reset); --
    end block;
    -- CP-element group 181:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	182 
    -- CP-element group 181: marked-predecessors 
    -- CP-element group 181: 	183 
    -- CP-element group 181: successors 
    -- CP-element group 181: 	183 
    -- CP-element group 181:  members (3) 
      -- CP-element group 181: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/WPIPE_d_out_buf_13022_update_start_
      -- CP-element group 181: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/WPIPE_d_out_buf_13022_Update/$entry
      -- CP-element group 181: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/WPIPE_d_out_buf_13022_Update/req
      -- 
    req_7325_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7325_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_6409_elements(181), ack => WPIPE_d_out_buf_13022_inst_req_1); -- 
    d_block_daemon_cp_element_group_181: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 2,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "d_block_daemon_cp_element_group_181"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= d_block_daemon_CP_6409_elements(182) & d_block_daemon_CP_6409_elements(183);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => d_block_daemon_CP_6409_elements(181), clk => clk, reset => reset); --
    end block;
    -- CP-element group 182:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	180 
    -- CP-element group 182: successors 
    -- CP-element group 182: 	181 
    -- CP-element group 182: marked-successors 
    -- CP-element group 182: 	177 
    -- CP-element group 182: 	180 
    -- CP-element group 182:  members (3) 
      -- CP-element group 182: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/WPIPE_d_out_buf_13022_sample_completed_
      -- CP-element group 182: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/WPIPE_d_out_buf_13022_Sample/$exit
      -- CP-element group 182: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/WPIPE_d_out_buf_13022_Sample/ack
      -- 
    ack_7321_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 182_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_d_out_buf_13022_inst_ack_0, ack => d_block_daemon_CP_6409_elements(182)); -- 
    -- CP-element group 183:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: 	181 
    -- CP-element group 183: successors 
    -- CP-element group 183: 	249 
    -- CP-element group 183: marked-successors 
    -- CP-element group 183: 	181 
    -- CP-element group 183:  members (3) 
      -- CP-element group 183: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/WPIPE_d_out_buf_13022_update_completed_
      -- CP-element group 183: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/WPIPE_d_out_buf_13022_Update/$exit
      -- CP-element group 183: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/WPIPE_d_out_buf_13022_Update/ack
      -- 
    ack_7326_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 183_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_d_out_buf_13022_inst_ack_1, ack => d_block_daemon_CP_6409_elements(183)); -- 
    -- CP-element group 184:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	63 
    -- CP-element group 184: marked-predecessors 
    -- CP-element group 184: 	186 
    -- CP-element group 184: successors 
    -- CP-element group 184: 	186 
    -- CP-element group 184:  members (3) 
      -- CP-element group 184: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/ADD_u15_u15_13028_sample_start_
      -- CP-element group 184: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/ADD_u15_u15_13028_Sample/$entry
      -- CP-element group 184: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/ADD_u15_u15_13028_Sample/rr
      -- 
    rr_7338_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7338_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_6409_elements(184), ack => ADD_u15_u15_13028_inst_req_0); -- 
    d_block_daemon_cp_element_group_184: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 2,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "d_block_daemon_cp_element_group_184"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= d_block_daemon_CP_6409_elements(63) & d_block_daemon_CP_6409_elements(186);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => d_block_daemon_CP_6409_elements(184), clk => clk, reset => reset); --
    end block;
    -- CP-element group 185:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	62 
    -- CP-element group 185: marked-predecessors 
    -- CP-element group 185: 	187 
    -- CP-element group 185: successors 
    -- CP-element group 185: 	187 
    -- CP-element group 185:  members (3) 
      -- CP-element group 185: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/ADD_u15_u15_13028_update_start_
      -- CP-element group 185: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/ADD_u15_u15_13028_Update/$entry
      -- CP-element group 185: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/ADD_u15_u15_13028_Update/cr
      -- 
    cr_7343_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7343_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_6409_elements(185), ack => ADD_u15_u15_13028_inst_req_1); -- 
    d_block_daemon_cp_element_group_185: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 2,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "d_block_daemon_cp_element_group_185"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= d_block_daemon_CP_6409_elements(62) & d_block_daemon_CP_6409_elements(187);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => d_block_daemon_CP_6409_elements(185), clk => clk, reset => reset); --
    end block;
    -- CP-element group 186:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	184 
    -- CP-element group 186: successors 
    -- CP-element group 186: marked-successors 
    -- CP-element group 186: 	61 
    -- CP-element group 186: 	184 
    -- CP-element group 186:  members (3) 
      -- CP-element group 186: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/ADD_u15_u15_13028_sample_completed_
      -- CP-element group 186: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/ADD_u15_u15_13028_Sample/$exit
      -- CP-element group 186: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/ADD_u15_u15_13028_Sample/ra
      -- 
    ra_7339_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 186_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u15_u15_13028_inst_ack_0, ack => d_block_daemon_CP_6409_elements(186)); -- 
    -- CP-element group 187:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: 	185 
    -- CP-element group 187: successors 
    -- CP-element group 187: 	188 
    -- CP-element group 187: marked-successors 
    -- CP-element group 187: 	60 
    -- CP-element group 187: 	185 
    -- CP-element group 187:  members (7) 
      -- CP-element group 187: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/ADD_u15_u15_13028_update_completed_
      -- CP-element group 187: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/ADD_u15_u15_13028_Update/$exit
      -- CP-element group 187: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/ADD_u15_u15_13028_Update/ca
      -- CP-element group 187: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_n_count_var_13031_sample_start_
      -- CP-element group 187: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_n_count_var_13031_sample_completed_
      -- CP-element group 187: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_n_count_var_13031_update_start_
      -- CP-element group 187: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/R_n_count_var_13031_update_completed_
      -- 
    ca_7344_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 187_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u15_u15_13028_inst_ack_1, ack => d_block_daemon_CP_6409_elements(187)); -- 
    -- CP-element group 188:  join  transition  bypass  pipeline-parent 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: 	187 
    -- CP-element group 188: 	58 
    -- CP-element group 188: successors 
    -- CP-element group 188: 	59 
    -- CP-element group 188:  members (12) 
      -- CP-element group 188: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/ULT_u15_u1_13033_sample_start_
      -- CP-element group 188: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/ULT_u15_u1_13033_sample_completed_
      -- CP-element group 188: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/ULT_u15_u1_13033_update_start_
      -- CP-element group 188: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/ULT_u15_u1_13033_update_completed_
      -- CP-element group 188: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/ULT_u15_u1_13033_Sample/$entry
      -- CP-element group 188: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/ULT_u15_u1_13033_Sample/$exit
      -- CP-element group 188: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/ULT_u15_u1_13033_Sample/rr
      -- CP-element group 188: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/ULT_u15_u1_13033_Sample/ra
      -- CP-element group 188: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/ULT_u15_u1_13033_Update/$entry
      -- CP-element group 188: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/ULT_u15_u1_13033_Update/$exit
      -- CP-element group 188: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/ULT_u15_u1_13033_Update/cr
      -- CP-element group 188: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/ULT_u15_u1_13033_Update/ca
      -- 
    d_block_daemon_cp_element_group_188: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 2,1 => 2);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "d_block_daemon_cp_element_group_188"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= d_block_daemon_CP_6409_elements(187) & d_block_daemon_CP_6409_elements(58);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => d_block_daemon_CP_6409_elements(188), clk => clk, reset => reset); --
    end block;
    -- CP-element group 189:  transition  bypass  pipeline-parent 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: 	54 
    -- CP-element group 189: successors 
    -- CP-element group 189: 	190 
    -- CP-element group 189:  members (1) 
      -- CP-element group 189: 	 branch_block_stmt_12832/do_while_stmt_12924/loop_exit/$entry
      -- 
    d_block_daemon_CP_6409_elements(189) <= d_block_daemon_CP_6409_elements(54);
    -- CP-element group 190:  transition  input  bypass  pipeline-parent 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: 	189 
    -- CP-element group 190: successors 
    -- CP-element group 190:  members (2) 
      -- CP-element group 190: 	 branch_block_stmt_12832/do_while_stmt_12924/loop_exit/$exit
      -- CP-element group 190: 	 branch_block_stmt_12832/do_while_stmt_12924/loop_exit/ack
      -- 
    ack_7370_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 190_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_12924_branch_ack_0, ack => d_block_daemon_CP_6409_elements(190)); -- 
    -- CP-element group 191:  transition  bypass  pipeline-parent 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: 	54 
    -- CP-element group 191: successors 
    -- CP-element group 191: 	192 
    -- CP-element group 191:  members (1) 
      -- CP-element group 191: 	 branch_block_stmt_12832/do_while_stmt_12924/loop_taken/$entry
      -- 
    d_block_daemon_CP_6409_elements(191) <= d_block_daemon_CP_6409_elements(54);
    -- CP-element group 192:  transition  input  bypass  pipeline-parent 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: 	191 
    -- CP-element group 192: successors 
    -- CP-element group 192:  members (2) 
      -- CP-element group 192: 	 branch_block_stmt_12832/do_while_stmt_12924/loop_taken/$exit
      -- CP-element group 192: 	 branch_block_stmt_12832/do_while_stmt_12924/loop_taken/ack
      -- 
    ack_7374_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 192_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_12924_branch_ack_1, ack => d_block_daemon_CP_6409_elements(192)); -- 
    -- CP-element group 193:  transition  bypass  pipeline-parent 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: 	52 
    -- CP-element group 193: successors 
    -- CP-element group 193: 	10 
    -- CP-element group 193:  members (1) 
      -- CP-element group 193: 	 branch_block_stmt_12832/do_while_stmt_12924/$exit
      -- 
    d_block_daemon_CP_6409_elements(193) <= d_block_daemon_CP_6409_elements(52);
    -- CP-element group 194:  transition  output  bypass 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: 	10 
    -- CP-element group 194: successors 
    -- CP-element group 194: 	195 
    -- CP-element group 194:  members (4) 
      -- CP-element group 194: 	 branch_block_stmt_12832/assign_stmt_13036/$entry
      -- CP-element group 194: 	 branch_block_stmt_12832/assign_stmt_13036/WPIPE_d_block_done_13034_sample_start_
      -- CP-element group 194: 	 branch_block_stmt_12832/assign_stmt_13036/WPIPE_d_block_done_13034_Sample/$entry
      -- CP-element group 194: 	 branch_block_stmt_12832/assign_stmt_13036/WPIPE_d_block_done_13034_Sample/req
      -- 
    req_7386_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7386_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_6409_elements(194), ack => WPIPE_d_block_done_13034_inst_req_0); -- 
    d_block_daemon_CP_6409_elements(194) <= d_block_daemon_CP_6409_elements(10);
    -- CP-element group 195:  transition  input  output  bypass 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: 	194 
    -- CP-element group 195: successors 
    -- CP-element group 195: 	196 
    -- CP-element group 195:  members (6) 
      -- CP-element group 195: 	 branch_block_stmt_12832/assign_stmt_13036/WPIPE_d_block_done_13034_sample_completed_
      -- CP-element group 195: 	 branch_block_stmt_12832/assign_stmt_13036/WPIPE_d_block_done_13034_update_start_
      -- CP-element group 195: 	 branch_block_stmt_12832/assign_stmt_13036/WPIPE_d_block_done_13034_Sample/$exit
      -- CP-element group 195: 	 branch_block_stmt_12832/assign_stmt_13036/WPIPE_d_block_done_13034_Sample/ack
      -- CP-element group 195: 	 branch_block_stmt_12832/assign_stmt_13036/WPIPE_d_block_done_13034_Update/$entry
      -- CP-element group 195: 	 branch_block_stmt_12832/assign_stmt_13036/WPIPE_d_block_done_13034_Update/req
      -- 
    ack_7387_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 195_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_d_block_done_13034_inst_ack_0, ack => d_block_daemon_CP_6409_elements(195)); -- 
    req_7391_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7391_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_6409_elements(195), ack => WPIPE_d_block_done_13034_inst_req_1); -- 
    -- CP-element group 196:  transition  input  bypass 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: 	195 
    -- CP-element group 196: successors 
    -- CP-element group 196: 	11 
    -- CP-element group 196:  members (4) 
      -- CP-element group 196: 	 branch_block_stmt_12832/assign_stmt_13036/$exit
      -- CP-element group 196: 	 branch_block_stmt_12832/assign_stmt_13036/WPIPE_d_block_done_13034_update_completed_
      -- CP-element group 196: 	 branch_block_stmt_12832/assign_stmt_13036/WPIPE_d_block_done_13034_Update/$exit
      -- CP-element group 196: 	 branch_block_stmt_12832/assign_stmt_13036/WPIPE_d_block_done_13034_Update/ack
      -- 
    ack_7392_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 196_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_d_block_done_13034_inst_ack_1, ack => d_block_daemon_CP_6409_elements(196)); -- 
    -- CP-element group 197:  transition  output  bypass 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: 	11 
    -- CP-element group 197: successors 
    -- CP-element group 197: 	198 
    -- CP-element group 197:  members (4) 
      -- CP-element group 197: 	 branch_block_stmt_12832/assign_stmt_13039/$entry
      -- CP-element group 197: 	 branch_block_stmt_12832/assign_stmt_13039/RPIPE_d_cmd_pipe_13038_sample_start_
      -- CP-element group 197: 	 branch_block_stmt_12832/assign_stmt_13039/RPIPE_d_cmd_pipe_13038_Sample/$entry
      -- CP-element group 197: 	 branch_block_stmt_12832/assign_stmt_13039/RPIPE_d_cmd_pipe_13038_Sample/rr
      -- 
    rr_7403_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7403_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_6409_elements(197), ack => RPIPE_d_cmd_pipe_13038_inst_req_0); -- 
    d_block_daemon_CP_6409_elements(197) <= d_block_daemon_CP_6409_elements(11);
    -- CP-element group 198:  transition  input  output  bypass 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: 	197 
    -- CP-element group 198: successors 
    -- CP-element group 198: 	199 
    -- CP-element group 198:  members (6) 
      -- CP-element group 198: 	 branch_block_stmt_12832/assign_stmt_13039/RPIPE_d_cmd_pipe_13038_sample_completed_
      -- CP-element group 198: 	 branch_block_stmt_12832/assign_stmt_13039/RPIPE_d_cmd_pipe_13038_update_start_
      -- CP-element group 198: 	 branch_block_stmt_12832/assign_stmt_13039/RPIPE_d_cmd_pipe_13038_Sample/$exit
      -- CP-element group 198: 	 branch_block_stmt_12832/assign_stmt_13039/RPIPE_d_cmd_pipe_13038_Sample/ra
      -- CP-element group 198: 	 branch_block_stmt_12832/assign_stmt_13039/RPIPE_d_cmd_pipe_13038_Update/$entry
      -- CP-element group 198: 	 branch_block_stmt_12832/assign_stmt_13039/RPIPE_d_cmd_pipe_13038_Update/cr
      -- 
    ra_7404_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 198_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_d_cmd_pipe_13038_inst_ack_0, ack => d_block_daemon_CP_6409_elements(198)); -- 
    cr_7408_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7408_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_6409_elements(198), ack => RPIPE_d_cmd_pipe_13038_inst_req_1); -- 
    -- CP-element group 199:  transition  input  bypass 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: 	198 
    -- CP-element group 199: successors 
    -- CP-element group 199: 	12 
    -- CP-element group 199:  members (4) 
      -- CP-element group 199: 	 branch_block_stmt_12832/assign_stmt_13039/$exit
      -- CP-element group 199: 	 branch_block_stmt_12832/assign_stmt_13039/RPIPE_d_cmd_pipe_13038_update_completed_
      -- CP-element group 199: 	 branch_block_stmt_12832/assign_stmt_13039/RPIPE_d_cmd_pipe_13038_Update/$exit
      -- CP-element group 199: 	 branch_block_stmt_12832/assign_stmt_13039/RPIPE_d_cmd_pipe_13038_Update/ca
      -- 
    ca_7409_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 199_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_d_cmd_pipe_13038_inst_ack_1, ack => d_block_daemon_CP_6409_elements(199)); -- 
    -- CP-element group 200:  join  fork  transition  bypass 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: 	12 
    -- CP-element group 200: successors 
    -- CP-element group 200: 	13 
    -- CP-element group 200:  members (50) 
      -- CP-element group 200: 	 branch_block_stmt_12832/assign_stmt_13043_to_assign_stmt_13051/R_d_new_cmd_13049_sample_start_
      -- CP-element group 200: 	 branch_block_stmt_12832/assign_stmt_13043_to_assign_stmt_13051/R_d_new_cmd_13049_update_start_
      -- CP-element group 200: 	 branch_block_stmt_12832/assign_stmt_13043_to_assign_stmt_13051/R_d_new_cmd_13049_sample_completed_
      -- CP-element group 200: 	 branch_block_stmt_12832/assign_stmt_13043_to_assign_stmt_13051/slice_13050_Update/ca
      -- CP-element group 200: 	 branch_block_stmt_12832/assign_stmt_13043_to_assign_stmt_13051/slice_13050_Update/cr
      -- CP-element group 200: 	 branch_block_stmt_12832/assign_stmt_13043_to_assign_stmt_13051/slice_13050_Update/$exit
      -- CP-element group 200: 	 branch_block_stmt_12832/assign_stmt_13043_to_assign_stmt_13051/slice_13050_Update/$entry
      -- CP-element group 200: 	 branch_block_stmt_12832/assign_stmt_13043_to_assign_stmt_13051/slice_13050_Sample/ra
      -- CP-element group 200: 	 branch_block_stmt_12832/assign_stmt_13043_to_assign_stmt_13051/slice_13050_Sample/rr
      -- CP-element group 200: 	 branch_block_stmt_12832/assign_stmt_13043_to_assign_stmt_13051/slice_13050_Sample/$exit
      -- CP-element group 200: 	 branch_block_stmt_12832/assign_stmt_13043_to_assign_stmt_13051/slice_13050_Sample/$entry
      -- CP-element group 200: 	 branch_block_stmt_12832/assign_stmt_13043_to_assign_stmt_13051/R_d_new_cmd_13049_update_completed_
      -- CP-element group 200: 	 branch_block_stmt_12832/assign_stmt_13043_to_assign_stmt_13051/$entry
      -- CP-element group 200: 	 branch_block_stmt_12832/assign_stmt_13043_to_assign_stmt_13051/$exit
      -- CP-element group 200: 	 branch_block_stmt_12832/assign_stmt_13043_to_assign_stmt_13051/slice_13042_sample_start_
      -- CP-element group 200: 	 branch_block_stmt_12832/assign_stmt_13043_to_assign_stmt_13051/slice_13042_sample_completed_
      -- CP-element group 200: 	 branch_block_stmt_12832/assign_stmt_13043_to_assign_stmt_13051/slice_13042_update_start_
      -- CP-element group 200: 	 branch_block_stmt_12832/assign_stmt_13043_to_assign_stmt_13051/slice_13042_update_completed_
      -- CP-element group 200: 	 branch_block_stmt_12832/assign_stmt_13043_to_assign_stmt_13051/R_d_new_cmd_13041_sample_start_
      -- CP-element group 200: 	 branch_block_stmt_12832/assign_stmt_13043_to_assign_stmt_13051/R_d_new_cmd_13041_sample_completed_
      -- CP-element group 200: 	 branch_block_stmt_12832/assign_stmt_13043_to_assign_stmt_13051/R_d_new_cmd_13041_update_start_
      -- CP-element group 200: 	 branch_block_stmt_12832/assign_stmt_13043_to_assign_stmt_13051/R_d_new_cmd_13041_update_completed_
      -- CP-element group 200: 	 branch_block_stmt_12832/assign_stmt_13043_to_assign_stmt_13051/slice_13042_Sample/$entry
      -- CP-element group 200: 	 branch_block_stmt_12832/assign_stmt_13043_to_assign_stmt_13051/slice_13042_Sample/$exit
      -- CP-element group 200: 	 branch_block_stmt_12832/assign_stmt_13043_to_assign_stmt_13051/slice_13042_Sample/rr
      -- CP-element group 200: 	 branch_block_stmt_12832/assign_stmt_13043_to_assign_stmt_13051/slice_13042_Sample/ra
      -- CP-element group 200: 	 branch_block_stmt_12832/assign_stmt_13043_to_assign_stmt_13051/slice_13042_Update/$entry
      -- CP-element group 200: 	 branch_block_stmt_12832/assign_stmt_13043_to_assign_stmt_13051/slice_13042_Update/$exit
      -- CP-element group 200: 	 branch_block_stmt_12832/assign_stmt_13043_to_assign_stmt_13051/slice_13042_Update/cr
      -- CP-element group 200: 	 branch_block_stmt_12832/assign_stmt_13043_to_assign_stmt_13051/slice_13042_Update/ca
      -- CP-element group 200: 	 branch_block_stmt_12832/assign_stmt_13043_to_assign_stmt_13051/slice_13046_sample_start_
      -- CP-element group 200: 	 branch_block_stmt_12832/assign_stmt_13043_to_assign_stmt_13051/slice_13046_sample_completed_
      -- CP-element group 200: 	 branch_block_stmt_12832/assign_stmt_13043_to_assign_stmt_13051/slice_13046_update_start_
      -- CP-element group 200: 	 branch_block_stmt_12832/assign_stmt_13043_to_assign_stmt_13051/slice_13046_update_completed_
      -- CP-element group 200: 	 branch_block_stmt_12832/assign_stmt_13043_to_assign_stmt_13051/R_d_new_cmd_13045_sample_start_
      -- CP-element group 200: 	 branch_block_stmt_12832/assign_stmt_13043_to_assign_stmt_13051/R_d_new_cmd_13045_sample_completed_
      -- CP-element group 200: 	 branch_block_stmt_12832/assign_stmt_13043_to_assign_stmt_13051/R_d_new_cmd_13045_update_start_
      -- CP-element group 200: 	 branch_block_stmt_12832/assign_stmt_13043_to_assign_stmt_13051/R_d_new_cmd_13045_update_completed_
      -- CP-element group 200: 	 branch_block_stmt_12832/assign_stmt_13043_to_assign_stmt_13051/slice_13046_Sample/$entry
      -- CP-element group 200: 	 branch_block_stmt_12832/assign_stmt_13043_to_assign_stmt_13051/slice_13046_Sample/$exit
      -- CP-element group 200: 	 branch_block_stmt_12832/assign_stmt_13043_to_assign_stmt_13051/slice_13046_Sample/rr
      -- CP-element group 200: 	 branch_block_stmt_12832/assign_stmt_13043_to_assign_stmt_13051/slice_13046_Sample/ra
      -- CP-element group 200: 	 branch_block_stmt_12832/assign_stmt_13043_to_assign_stmt_13051/slice_13046_Update/$entry
      -- CP-element group 200: 	 branch_block_stmt_12832/assign_stmt_13043_to_assign_stmt_13051/slice_13046_Update/$exit
      -- CP-element group 200: 	 branch_block_stmt_12832/assign_stmt_13043_to_assign_stmt_13051/slice_13046_Update/cr
      -- CP-element group 200: 	 branch_block_stmt_12832/assign_stmt_13043_to_assign_stmt_13051/slice_13046_Update/ca
      -- CP-element group 200: 	 branch_block_stmt_12832/assign_stmt_13043_to_assign_stmt_13051/slice_13050_sample_start_
      -- CP-element group 200: 	 branch_block_stmt_12832/assign_stmt_13043_to_assign_stmt_13051/slice_13050_sample_completed_
      -- CP-element group 200: 	 branch_block_stmt_12832/assign_stmt_13043_to_assign_stmt_13051/slice_13050_update_start_
      -- CP-element group 200: 	 branch_block_stmt_12832/assign_stmt_13043_to_assign_stmt_13051/slice_13050_update_completed_
      -- 
    d_block_daemon_CP_6409_elements(200) <= d_block_daemon_CP_6409_elements(12);
    -- CP-element group 201:  transition  bypass 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: 	13 
    -- CP-element group 201: successors 
    -- CP-element group 201:  members (1) 
      -- CP-element group 201: 	 branch_block_stmt_12832/if_stmt_13052_dead_link/$entry
      -- 
    d_block_daemon_CP_6409_elements(201) <= d_block_daemon_CP_6409_elements(13);
    -- CP-element group 202:  transition  output  bypass 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: 	13 
    -- CP-element group 202: successors 
    -- CP-element group 202: 	203 
    -- CP-element group 202:  members (17) 
      -- CP-element group 202: 	 branch_block_stmt_12832/if_stmt_13052_eval_test/EQ_u1_u1_13055/SplitProtocol/Sample/rr
      -- CP-element group 202: 	 branch_block_stmt_12832/if_stmt_13052_eval_test/EQ_u1_u1_13055/SplitProtocol/Sample/$exit
      -- CP-element group 202: 	 branch_block_stmt_12832/if_stmt_13052_eval_test/EQ_u1_u1_13055/SplitProtocol/Sample/$entry
      -- CP-element group 202: 	 branch_block_stmt_12832/if_stmt_13052_eval_test/EQ_u1_u1_13055/SplitProtocol/$exit
      -- CP-element group 202: 	 branch_block_stmt_12832/if_stmt_13052_eval_test/EQ_u1_u1_13055/SplitProtocol/$entry
      -- CP-element group 202: 	 branch_block_stmt_12832/if_stmt_13052_eval_test/EQ_u1_u1_13055/EQ_u1_u1_13055_inputs/$exit
      -- CP-element group 202: 	 branch_block_stmt_12832/if_stmt_13052_eval_test/EQ_u1_u1_13055/EQ_u1_u1_13055_inputs/$entry
      -- CP-element group 202: 	 branch_block_stmt_12832/if_stmt_13052_eval_test/EQ_u1_u1_13055/$exit
      -- CP-element group 202: 	 branch_block_stmt_12832/if_stmt_13052_eval_test/EQ_u1_u1_13055/$entry
      -- CP-element group 202: 	 branch_block_stmt_12832/if_stmt_13052_eval_test/$exit
      -- CP-element group 202: 	 branch_block_stmt_12832/if_stmt_13052_eval_test/$entry
      -- CP-element group 202: 	 branch_block_stmt_12832/if_stmt_13052_eval_test/branch_req
      -- CP-element group 202: 	 branch_block_stmt_12832/if_stmt_13052_eval_test/EQ_u1_u1_13055/SplitProtocol/Update/ca
      -- CP-element group 202: 	 branch_block_stmt_12832/if_stmt_13052_eval_test/EQ_u1_u1_13055/SplitProtocol/Update/cr
      -- CP-element group 202: 	 branch_block_stmt_12832/if_stmt_13052_eval_test/EQ_u1_u1_13055/SplitProtocol/Update/$exit
      -- CP-element group 202: 	 branch_block_stmt_12832/if_stmt_13052_eval_test/EQ_u1_u1_13055/SplitProtocol/Update/$entry
      -- CP-element group 202: 	 branch_block_stmt_12832/if_stmt_13052_eval_test/EQ_u1_u1_13055/SplitProtocol/Sample/ra
      -- 
    branch_req_7493_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_7493_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_6409_elements(202), ack => if_stmt_13052_branch_req_0); -- 
    d_block_daemon_CP_6409_elements(202) <= d_block_daemon_CP_6409_elements(13);
    -- CP-element group 203:  branch  place  bypass 
    -- CP-element group 203: predecessors 
    -- CP-element group 203: 	202 
    -- CP-element group 203: successors 
    -- CP-element group 203: 	206 
    -- CP-element group 203: 	204 
    -- CP-element group 203:  members (1) 
      -- CP-element group 203: 	 branch_block_stmt_12832/EQ_u1_u1_13055_place
      -- 
    d_block_daemon_CP_6409_elements(203) <= d_block_daemon_CP_6409_elements(202);
    -- CP-element group 204:  transition  bypass 
    -- CP-element group 204: predecessors 
    -- CP-element group 204: 	203 
    -- CP-element group 204: successors 
    -- CP-element group 204: 	205 
    -- CP-element group 204:  members (1) 
      -- CP-element group 204: 	 branch_block_stmt_12832/if_stmt_13052_if_link/$entry
      -- 
    d_block_daemon_CP_6409_elements(204) <= d_block_daemon_CP_6409_elements(203);
    -- CP-element group 205:  transition  input  bypass 
    -- CP-element group 205: predecessors 
    -- CP-element group 205: 	204 
    -- CP-element group 205: successors 
    -- CP-element group 205: 	208 
    -- CP-element group 205:  members (2) 
      -- CP-element group 205: 	 branch_block_stmt_12832/if_stmt_13052_if_link/if_choice_transition
      -- CP-element group 205: 	 branch_block_stmt_12832/if_stmt_13052_if_link/$exit
      -- 
    if_choice_transition_7498_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 205_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_13052_branch_ack_1, ack => d_block_daemon_CP_6409_elements(205)); -- 
    -- CP-element group 206:  transition  bypass 
    -- CP-element group 206: predecessors 
    -- CP-element group 206: 	203 
    -- CP-element group 206: successors 
    -- CP-element group 206: 	207 
    -- CP-element group 206:  members (1) 
      -- CP-element group 206: 	 branch_block_stmt_12832/if_stmt_13052_else_link/$entry
      -- 
    d_block_daemon_CP_6409_elements(206) <= d_block_daemon_CP_6409_elements(203);
    -- CP-element group 207:  transition  input  bypass 
    -- CP-element group 207: predecessors 
    -- CP-element group 207: 	206 
    -- CP-element group 207: successors 
    -- CP-element group 207: 	209 
    -- CP-element group 207:  members (2) 
      -- CP-element group 207: 	 branch_block_stmt_12832/if_stmt_13052_else_link/else_choice_transition
      -- CP-element group 207: 	 branch_block_stmt_12832/if_stmt_13052_else_link/$exit
      -- 
    else_choice_transition_7502_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 207_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_13052_branch_ack_0, ack => d_block_daemon_CP_6409_elements(207)); -- 
    -- CP-element group 208:  place  bypass 
    -- CP-element group 208: predecessors 
    -- CP-element group 208: 	205 
    -- CP-element group 208: successors 
    -- CP-element group 208: 	224 
    -- CP-element group 208:  members (1) 
      -- CP-element group 208: 	 branch_block_stmt_12832/GotNewKey
      -- 
    d_block_daemon_CP_6409_elements(208) <= d_block_daemon_CP_6409_elements(205);
    -- CP-element group 209:  place  bypass 
    -- CP-element group 209: predecessors 
    -- CP-element group 209: 	207 
    -- CP-element group 209: successors 
    -- CP-element group 209: 	242 
    -- CP-element group 209:  members (1) 
      -- CP-element group 209: 	 branch_block_stmt_12832/NotGotNewKey
      -- 
    d_block_daemon_CP_6409_elements(209) <= d_block_daemon_CP_6409_elements(207);
    -- CP-element group 210:  transition  bypass 
    -- CP-element group 210: predecessors 
    -- CP-element group 210: 	2 
    -- CP-element group 210: successors 
    -- CP-element group 210:  members (1) 
      -- CP-element group 210: 	 branch_block_stmt_12832/merge_stmt_12836_dead_link/$entry
      -- 
    d_block_daemon_CP_6409_elements(210) <= d_block_daemon_CP_6409_elements(2);
    -- CP-element group 211:  transition  bypass 
    -- CP-element group 211: predecessors 
    -- CP-element group 211: 	2 
    -- CP-element group 211: successors 
    -- CP-element group 211: 	213 
    -- CP-element group 211:  members (2) 
      -- CP-element group 211: 	 branch_block_stmt_12832/merge_stmt_12836__entry___PhiReq/$exit
      -- CP-element group 211: 	 branch_block_stmt_12832/merge_stmt_12836__entry___PhiReq/$entry
      -- 
    d_block_daemon_CP_6409_elements(211) <= d_block_daemon_CP_6409_elements(2);
    -- CP-element group 212:  transition  bypass 
    -- CP-element group 212: predecessors 
    -- CP-element group 212: 	28 
    -- CP-element group 212: successors 
    -- CP-element group 212: 	213 
    -- CP-element group 212:  members (2) 
      -- CP-element group 212: 	 branch_block_stmt_12832/NotGotCmd_PhiReq/$exit
      -- CP-element group 212: 	 branch_block_stmt_12832/NotGotCmd_PhiReq/$entry
      -- 
    d_block_daemon_CP_6409_elements(212) <= d_block_daemon_CP_6409_elements(28);
    -- CP-element group 213:  merge  place  bypass 
    -- CP-element group 213: predecessors 
    -- CP-element group 213: 	211 
    -- CP-element group 213: 	212 
    -- CP-element group 213: successors 
    -- CP-element group 213: 	214 
    -- CP-element group 213:  members (1) 
      -- CP-element group 213: 	 branch_block_stmt_12832/merge_stmt_12836_PhiReqMerge
      -- 
    d_block_daemon_CP_6409_elements(213) <= OrReduce(d_block_daemon_CP_6409_elements(211) & d_block_daemon_CP_6409_elements(212));
    -- CP-element group 214:  transition  bypass 
    -- CP-element group 214: predecessors 
    -- CP-element group 214: 	213 
    -- CP-element group 214: successors 
    -- CP-element group 214: 	3 
    -- CP-element group 214:  members (3) 
      -- CP-element group 214: 	 branch_block_stmt_12832/merge_stmt_12836_PhiAck/$entry
      -- CP-element group 214: 	 branch_block_stmt_12832/merge_stmt_12836_PhiAck/$exit
      -- CP-element group 214: 	 branch_block_stmt_12832/merge_stmt_12836_PhiAck/dummy
      -- 
    d_block_daemon_CP_6409_elements(214) <= d_block_daemon_CP_6409_elements(213);
    -- CP-element group 215:  transition  bypass 
    -- CP-element group 215: predecessors 
    -- CP-element group 215: 	6 
    -- CP-element group 215: successors 
    -- CP-element group 215:  members (1) 
      -- CP-element group 215: 	 branch_block_stmt_12832/merge_stmt_12858_dead_link/$entry
      -- 
    d_block_daemon_CP_6409_elements(215) <= d_block_daemon_CP_6409_elements(6);
    -- CP-element group 216:  fork  transition  output  bypass 
    -- CP-element group 216: predecessors 
    -- CP-element group 216: 	6 
    -- CP-element group 216: successors 
    -- CP-element group 216: 	217 
    -- CP-element group 216: 	218 
    -- CP-element group 216: 	220 
    -- CP-element group 216: 	221 
    -- CP-element group 216:  members (15) 
      -- CP-element group 216: 	 branch_block_stmt_12832/merge_stmt_12858__entry___PhiReq/$entry
      -- CP-element group 216: 	 branch_block_stmt_12832/merge_stmt_12858__entry___PhiReq/phi_stmt_12859/phi_stmt_12859_sources/$entry
      -- CP-element group 216: 	 branch_block_stmt_12832/merge_stmt_12858__entry___PhiReq/phi_stmt_12863/phi_stmt_12863_sources/$entry
      -- CP-element group 216: 	 branch_block_stmt_12832/merge_stmt_12858__entry___PhiReq/phi_stmt_12863/$entry
      -- CP-element group 216: 	 branch_block_stmt_12832/merge_stmt_12858__entry___PhiReq/phi_stmt_12859/$entry
      -- CP-element group 216: 	 branch_block_stmt_12832/merge_stmt_12858__entry___PhiReq/phi_stmt_12859/phi_stmt_12859_sources/Interlock/Update/req
      -- CP-element group 216: 	 branch_block_stmt_12832/merge_stmt_12858__entry___PhiReq/phi_stmt_12859/phi_stmt_12859_sources/Interlock/Update/$entry
      -- CP-element group 216: 	 branch_block_stmt_12832/merge_stmt_12858__entry___PhiReq/phi_stmt_12859/phi_stmt_12859_sources/Interlock/Sample/req
      -- CP-element group 216: 	 branch_block_stmt_12832/merge_stmt_12858__entry___PhiReq/phi_stmt_12863/phi_stmt_12863_sources/Interlock/Update/req
      -- CP-element group 216: 	 branch_block_stmt_12832/merge_stmt_12858__entry___PhiReq/phi_stmt_12859/phi_stmt_12859_sources/Interlock/Sample/$entry
      -- CP-element group 216: 	 branch_block_stmt_12832/merge_stmt_12858__entry___PhiReq/phi_stmt_12863/phi_stmt_12863_sources/Interlock/Update/$entry
      -- CP-element group 216: 	 branch_block_stmt_12832/merge_stmt_12858__entry___PhiReq/phi_stmt_12859/phi_stmt_12859_sources/Interlock/$entry
      -- CP-element group 216: 	 branch_block_stmt_12832/merge_stmt_12858__entry___PhiReq/phi_stmt_12863/phi_stmt_12863_sources/Interlock/Sample/req
      -- CP-element group 216: 	 branch_block_stmt_12832/merge_stmt_12858__entry___PhiReq/phi_stmt_12863/phi_stmt_12863_sources/Interlock/Sample/$entry
      -- CP-element group 216: 	 branch_block_stmt_12832/merge_stmt_12858__entry___PhiReq/phi_stmt_12863/phi_stmt_12863_sources/Interlock/$entry
      -- 
    req_7539_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7539_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_6409_elements(216), ack => d_init_key_12851_12861_buf_req_0); -- 
    req_7544_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7544_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_6409_elements(216), ack => d_init_key_12851_12861_buf_req_1); -- 
    req_7559_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7559_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_6409_elements(216), ack => d_init_count_12847_12865_buf_req_0); -- 
    req_7564_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7564_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_6409_elements(216), ack => d_init_count_12847_12865_buf_req_1); -- 
    d_block_daemon_CP_6409_elements(216) <= d_block_daemon_CP_6409_elements(6);
    -- CP-element group 217:  transition  input  bypass 
    -- CP-element group 217: predecessors 
    -- CP-element group 217: 	216 
    -- CP-element group 217: successors 
    -- CP-element group 217: 	219 
    -- CP-element group 217:  members (2) 
      -- CP-element group 217: 	 branch_block_stmt_12832/merge_stmt_12858__entry___PhiReq/phi_stmt_12859/phi_stmt_12859_sources/Interlock/Sample/ack
      -- CP-element group 217: 	 branch_block_stmt_12832/merge_stmt_12858__entry___PhiReq/phi_stmt_12859/phi_stmt_12859_sources/Interlock/Sample/$exit
      -- 
    ack_7540_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 217_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_init_key_12851_12861_buf_ack_0, ack => d_block_daemon_CP_6409_elements(217)); -- 
    -- CP-element group 218:  transition  input  bypass 
    -- CP-element group 218: predecessors 
    -- CP-element group 218: 	216 
    -- CP-element group 218: successors 
    -- CP-element group 218: 	219 
    -- CP-element group 218:  members (2) 
      -- CP-element group 218: 	 branch_block_stmt_12832/merge_stmt_12858__entry___PhiReq/phi_stmt_12859/phi_stmt_12859_sources/Interlock/Update/ack
      -- CP-element group 218: 	 branch_block_stmt_12832/merge_stmt_12858__entry___PhiReq/phi_stmt_12859/phi_stmt_12859_sources/Interlock/Update/$exit
      -- 
    ack_7545_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 218_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_init_key_12851_12861_buf_ack_1, ack => d_block_daemon_CP_6409_elements(218)); -- 
    -- CP-element group 219:  join  transition  output  bypass 
    -- CP-element group 219: predecessors 
    -- CP-element group 219: 	217 
    -- CP-element group 219: 	218 
    -- CP-element group 219: successors 
    -- CP-element group 219: 	223 
    -- CP-element group 219:  members (4) 
      -- CP-element group 219: 	 branch_block_stmt_12832/merge_stmt_12858__entry___PhiReq/phi_stmt_12859/phi_stmt_12859_sources/$exit
      -- CP-element group 219: 	 branch_block_stmt_12832/merge_stmt_12858__entry___PhiReq/phi_stmt_12859/$exit
      -- CP-element group 219: 	 branch_block_stmt_12832/merge_stmt_12858__entry___PhiReq/phi_stmt_12859/phi_stmt_12859_req
      -- CP-element group 219: 	 branch_block_stmt_12832/merge_stmt_12858__entry___PhiReq/phi_stmt_12859/phi_stmt_12859_sources/Interlock/$exit
      -- 
    phi_stmt_12859_req_7546_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_12859_req_7546_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_6409_elements(219), ack => phi_stmt_12859_req_0); -- 
    d_block_daemon_cp_element_group_219: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "d_block_daemon_cp_element_group_219"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= d_block_daemon_CP_6409_elements(217) & d_block_daemon_CP_6409_elements(218);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => d_block_daemon_CP_6409_elements(219), clk => clk, reset => reset); --
    end block;
    -- CP-element group 220:  transition  input  bypass 
    -- CP-element group 220: predecessors 
    -- CP-element group 220: 	216 
    -- CP-element group 220: successors 
    -- CP-element group 220: 	222 
    -- CP-element group 220:  members (2) 
      -- CP-element group 220: 	 branch_block_stmt_12832/merge_stmt_12858__entry___PhiReq/phi_stmt_12863/phi_stmt_12863_sources/Interlock/Sample/ack
      -- CP-element group 220: 	 branch_block_stmt_12832/merge_stmt_12858__entry___PhiReq/phi_stmt_12863/phi_stmt_12863_sources/Interlock/Sample/$exit
      -- 
    ack_7560_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 220_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_init_count_12847_12865_buf_ack_0, ack => d_block_daemon_CP_6409_elements(220)); -- 
    -- CP-element group 221:  transition  input  bypass 
    -- CP-element group 221: predecessors 
    -- CP-element group 221: 	216 
    -- CP-element group 221: successors 
    -- CP-element group 221: 	222 
    -- CP-element group 221:  members (2) 
      -- CP-element group 221: 	 branch_block_stmt_12832/merge_stmt_12858__entry___PhiReq/phi_stmt_12863/phi_stmt_12863_sources/Interlock/Update/ack
      -- CP-element group 221: 	 branch_block_stmt_12832/merge_stmt_12858__entry___PhiReq/phi_stmt_12863/phi_stmt_12863_sources/Interlock/Update/$exit
      -- 
    ack_7565_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 221_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_init_count_12847_12865_buf_ack_1, ack => d_block_daemon_CP_6409_elements(221)); -- 
    -- CP-element group 222:  join  transition  output  bypass 
    -- CP-element group 222: predecessors 
    -- CP-element group 222: 	220 
    -- CP-element group 222: 	221 
    -- CP-element group 222: successors 
    -- CP-element group 222: 	223 
    -- CP-element group 222:  members (4) 
      -- CP-element group 222: 	 branch_block_stmt_12832/merge_stmt_12858__entry___PhiReq/phi_stmt_12863/phi_stmt_12863_sources/$exit
      -- CP-element group 222: 	 branch_block_stmt_12832/merge_stmt_12858__entry___PhiReq/phi_stmt_12863/$exit
      -- CP-element group 222: 	 branch_block_stmt_12832/merge_stmt_12858__entry___PhiReq/phi_stmt_12863/phi_stmt_12863_req
      -- CP-element group 222: 	 branch_block_stmt_12832/merge_stmt_12858__entry___PhiReq/phi_stmt_12863/phi_stmt_12863_sources/Interlock/$exit
      -- 
    phi_stmt_12863_req_7566_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_12863_req_7566_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_6409_elements(222), ack => phi_stmt_12863_req_0); -- 
    d_block_daemon_cp_element_group_222: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "d_block_daemon_cp_element_group_222"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= d_block_daemon_CP_6409_elements(220) & d_block_daemon_CP_6409_elements(221);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => d_block_daemon_CP_6409_elements(222), clk => clk, reset => reset); --
    end block;
    -- CP-element group 223:  join  transition  bypass 
    -- CP-element group 223: predecessors 
    -- CP-element group 223: 	219 
    -- CP-element group 223: 	222 
    -- CP-element group 223: successors 
    -- CP-element group 223: 	232 
    -- CP-element group 223:  members (1) 
      -- CP-element group 223: 	 branch_block_stmt_12832/merge_stmt_12858__entry___PhiReq/$exit
      -- 
    d_block_daemon_cp_element_group_223: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "d_block_daemon_cp_element_group_223"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= d_block_daemon_CP_6409_elements(219) & d_block_daemon_CP_6409_elements(222);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => d_block_daemon_CP_6409_elements(223), clk => clk, reset => reset); --
    end block;
    -- CP-element group 224:  fork  transition  output  bypass 
    -- CP-element group 224: predecessors 
    -- CP-element group 224: 	208 
    -- CP-element group 224: successors 
    -- CP-element group 224: 	225 
    -- CP-element group 224: 	226 
    -- CP-element group 224: 	228 
    -- CP-element group 224: 	229 
    -- CP-element group 224:  members (15) 
      -- CP-element group 224: 	 branch_block_stmt_12832/GotNewKey_PhiReq/phi_stmt_12863/phi_stmt_12863_sources/Interlock/$entry
      -- CP-element group 224: 	 branch_block_stmt_12832/GotNewKey_PhiReq/phi_stmt_12859/phi_stmt_12859_sources/Interlock/Sample/$entry
      -- CP-element group 224: 	 branch_block_stmt_12832/GotNewKey_PhiReq/phi_stmt_12859/phi_stmt_12859_sources/Interlock/$entry
      -- CP-element group 224: 	 branch_block_stmt_12832/GotNewKey_PhiReq/phi_stmt_12863/phi_stmt_12863_sources/$entry
      -- CP-element group 224: 	 branch_block_stmt_12832/GotNewKey_PhiReq/phi_stmt_12859/phi_stmt_12859_sources/$entry
      -- CP-element group 224: 	 branch_block_stmt_12832/GotNewKey_PhiReq/phi_stmt_12859/$entry
      -- CP-element group 224: 	 branch_block_stmt_12832/GotNewKey_PhiReq/$entry
      -- CP-element group 224: 	 branch_block_stmt_12832/GotNewKey_PhiReq/phi_stmt_12863/$entry
      -- CP-element group 224: 	 branch_block_stmt_12832/GotNewKey_PhiReq/phi_stmt_12863/phi_stmt_12863_sources/Interlock/Update/req
      -- CP-element group 224: 	 branch_block_stmt_12832/GotNewKey_PhiReq/phi_stmt_12859/phi_stmt_12859_sources/Interlock/Update/req
      -- CP-element group 224: 	 branch_block_stmt_12832/GotNewKey_PhiReq/phi_stmt_12863/phi_stmt_12863_sources/Interlock/Update/$entry
      -- CP-element group 224: 	 branch_block_stmt_12832/GotNewKey_PhiReq/phi_stmt_12859/phi_stmt_12859_sources/Interlock/Update/$entry
      -- CP-element group 224: 	 branch_block_stmt_12832/GotNewKey_PhiReq/phi_stmt_12863/phi_stmt_12863_sources/Interlock/Sample/req
      -- CP-element group 224: 	 branch_block_stmt_12832/GotNewKey_PhiReq/phi_stmt_12863/phi_stmt_12863_sources/Interlock/Sample/$entry
      -- CP-element group 224: 	 branch_block_stmt_12832/GotNewKey_PhiReq/phi_stmt_12859/phi_stmt_12859_sources/Interlock/Sample/req
      -- 
    req_7582_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7582_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_6409_elements(224), ack => d_new_key_13051_12862_buf_req_0); -- 
    req_7587_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7587_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_6409_elements(224), ack => d_new_key_13051_12862_buf_req_1); -- 
    req_7602_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7602_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_6409_elements(224), ack => d_new_count_13047_12866_buf_req_0); -- 
    req_7607_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7607_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_6409_elements(224), ack => d_new_count_13047_12866_buf_req_1); -- 
    d_block_daemon_CP_6409_elements(224) <= d_block_daemon_CP_6409_elements(208);
    -- CP-element group 225:  transition  input  bypass 
    -- CP-element group 225: predecessors 
    -- CP-element group 225: 	224 
    -- CP-element group 225: successors 
    -- CP-element group 225: 	227 
    -- CP-element group 225:  members (2) 
      -- CP-element group 225: 	 branch_block_stmt_12832/GotNewKey_PhiReq/phi_stmt_12859/phi_stmt_12859_sources/Interlock/Sample/$exit
      -- CP-element group 225: 	 branch_block_stmt_12832/GotNewKey_PhiReq/phi_stmt_12859/phi_stmt_12859_sources/Interlock/Sample/ack
      -- 
    ack_7583_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 225_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_new_key_13051_12862_buf_ack_0, ack => d_block_daemon_CP_6409_elements(225)); -- 
    -- CP-element group 226:  transition  input  bypass 
    -- CP-element group 226: predecessors 
    -- CP-element group 226: 	224 
    -- CP-element group 226: successors 
    -- CP-element group 226: 	227 
    -- CP-element group 226:  members (2) 
      -- CP-element group 226: 	 branch_block_stmt_12832/GotNewKey_PhiReq/phi_stmt_12859/phi_stmt_12859_sources/Interlock/Update/ack
      -- CP-element group 226: 	 branch_block_stmt_12832/GotNewKey_PhiReq/phi_stmt_12859/phi_stmt_12859_sources/Interlock/Update/$exit
      -- 
    ack_7588_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 226_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_new_key_13051_12862_buf_ack_1, ack => d_block_daemon_CP_6409_elements(226)); -- 
    -- CP-element group 227:  join  transition  output  bypass 
    -- CP-element group 227: predecessors 
    -- CP-element group 227: 	225 
    -- CP-element group 227: 	226 
    -- CP-element group 227: successors 
    -- CP-element group 227: 	231 
    -- CP-element group 227:  members (4) 
      -- CP-element group 227: 	 branch_block_stmt_12832/GotNewKey_PhiReq/phi_stmt_12859/phi_stmt_12859_sources/Interlock/$exit
      -- CP-element group 227: 	 branch_block_stmt_12832/GotNewKey_PhiReq/phi_stmt_12859/phi_stmt_12859_sources/$exit
      -- CP-element group 227: 	 branch_block_stmt_12832/GotNewKey_PhiReq/phi_stmt_12859/$exit
      -- CP-element group 227: 	 branch_block_stmt_12832/GotNewKey_PhiReq/phi_stmt_12859/phi_stmt_12859_req
      -- 
    phi_stmt_12859_req_7589_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_12859_req_7589_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_6409_elements(227), ack => phi_stmt_12859_req_1); -- 
    d_block_daemon_cp_element_group_227: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "d_block_daemon_cp_element_group_227"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= d_block_daemon_CP_6409_elements(225) & d_block_daemon_CP_6409_elements(226);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => d_block_daemon_CP_6409_elements(227), clk => clk, reset => reset); --
    end block;
    -- CP-element group 228:  transition  input  bypass 
    -- CP-element group 228: predecessors 
    -- CP-element group 228: 	224 
    -- CP-element group 228: successors 
    -- CP-element group 228: 	230 
    -- CP-element group 228:  members (2) 
      -- CP-element group 228: 	 branch_block_stmt_12832/GotNewKey_PhiReq/phi_stmt_12863/phi_stmt_12863_sources/Interlock/Sample/ack
      -- CP-element group 228: 	 branch_block_stmt_12832/GotNewKey_PhiReq/phi_stmt_12863/phi_stmt_12863_sources/Interlock/Sample/$exit
      -- 
    ack_7603_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 228_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_new_count_13047_12866_buf_ack_0, ack => d_block_daemon_CP_6409_elements(228)); -- 
    -- CP-element group 229:  transition  input  bypass 
    -- CP-element group 229: predecessors 
    -- CP-element group 229: 	224 
    -- CP-element group 229: successors 
    -- CP-element group 229: 	230 
    -- CP-element group 229:  members (2) 
      -- CP-element group 229: 	 branch_block_stmt_12832/GotNewKey_PhiReq/phi_stmt_12863/phi_stmt_12863_sources/Interlock/Update/ack
      -- CP-element group 229: 	 branch_block_stmt_12832/GotNewKey_PhiReq/phi_stmt_12863/phi_stmt_12863_sources/Interlock/Update/$exit
      -- 
    ack_7608_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 229_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_new_count_13047_12866_buf_ack_1, ack => d_block_daemon_CP_6409_elements(229)); -- 
    -- CP-element group 230:  join  transition  output  bypass 
    -- CP-element group 230: predecessors 
    -- CP-element group 230: 	228 
    -- CP-element group 230: 	229 
    -- CP-element group 230: successors 
    -- CP-element group 230: 	231 
    -- CP-element group 230:  members (4) 
      -- CP-element group 230: 	 branch_block_stmt_12832/GotNewKey_PhiReq/phi_stmt_12863/phi_stmt_12863_sources/Interlock/$exit
      -- CP-element group 230: 	 branch_block_stmt_12832/GotNewKey_PhiReq/phi_stmt_12863/phi_stmt_12863_req
      -- CP-element group 230: 	 branch_block_stmt_12832/GotNewKey_PhiReq/phi_stmt_12863/phi_stmt_12863_sources/$exit
      -- CP-element group 230: 	 branch_block_stmt_12832/GotNewKey_PhiReq/phi_stmt_12863/$exit
      -- 
    phi_stmt_12863_req_7609_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_12863_req_7609_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_6409_elements(230), ack => phi_stmt_12863_req_1); -- 
    d_block_daemon_cp_element_group_230: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "d_block_daemon_cp_element_group_230"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= d_block_daemon_CP_6409_elements(228) & d_block_daemon_CP_6409_elements(229);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => d_block_daemon_CP_6409_elements(230), clk => clk, reset => reset); --
    end block;
    -- CP-element group 231:  join  transition  bypass 
    -- CP-element group 231: predecessors 
    -- CP-element group 231: 	227 
    -- CP-element group 231: 	230 
    -- CP-element group 231: successors 
    -- CP-element group 231: 	232 
    -- CP-element group 231:  members (1) 
      -- CP-element group 231: 	 branch_block_stmt_12832/GotNewKey_PhiReq/$exit
      -- 
    d_block_daemon_cp_element_group_231: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "d_block_daemon_cp_element_group_231"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= d_block_daemon_CP_6409_elements(227) & d_block_daemon_CP_6409_elements(230);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => d_block_daemon_CP_6409_elements(231), clk => clk, reset => reset); --
    end block;
    -- CP-element group 232:  merge  place  bypass 
    -- CP-element group 232: predecessors 
    -- CP-element group 232: 	223 
    -- CP-element group 232: 	231 
    -- CP-element group 232: successors 
    -- CP-element group 232: 	233 
    -- CP-element group 232:  members (1) 
      -- CP-element group 232: 	 branch_block_stmt_12832/merge_stmt_12858_PhiReqMerge
      -- 
    d_block_daemon_CP_6409_elements(232) <= OrReduce(d_block_daemon_CP_6409_elements(223) & d_block_daemon_CP_6409_elements(231));
    -- CP-element group 233:  fork  transition  bypass 
    -- CP-element group 233: predecessors 
    -- CP-element group 233: 	232 
    -- CP-element group 233: successors 
    -- CP-element group 233: 	234 
    -- CP-element group 233: 	235 
    -- CP-element group 233:  members (1) 
      -- CP-element group 233: 	 branch_block_stmt_12832/merge_stmt_12858_PhiAck/$entry
      -- 
    d_block_daemon_CP_6409_elements(233) <= d_block_daemon_CP_6409_elements(232);
    -- CP-element group 234:  transition  input  bypass 
    -- CP-element group 234: predecessors 
    -- CP-element group 234: 	233 
    -- CP-element group 234: successors 
    -- CP-element group 234: 	236 
    -- CP-element group 234:  members (1) 
      -- CP-element group 234: 	 branch_block_stmt_12832/merge_stmt_12858_PhiAck/phi_stmt_12859_ack
      -- 
    phi_stmt_12859_ack_7614_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 234_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_12859_ack_0, ack => d_block_daemon_CP_6409_elements(234)); -- 
    -- CP-element group 235:  transition  input  bypass 
    -- CP-element group 235: predecessors 
    -- CP-element group 235: 	233 
    -- CP-element group 235: successors 
    -- CP-element group 235: 	236 
    -- CP-element group 235:  members (1) 
      -- CP-element group 235: 	 branch_block_stmt_12832/merge_stmt_12858_PhiAck/phi_stmt_12863_ack
      -- 
    phi_stmt_12863_ack_7615_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 235_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_12863_ack_0, ack => d_block_daemon_CP_6409_elements(235)); -- 
    -- CP-element group 236:  join  transition  bypass 
    -- CP-element group 236: predecessors 
    -- CP-element group 236: 	234 
    -- CP-element group 236: 	235 
    -- CP-element group 236: successors 
    -- CP-element group 236: 	7 
    -- CP-element group 236:  members (1) 
      -- CP-element group 236: 	 branch_block_stmt_12832/merge_stmt_12858_PhiAck/$exit
      -- 
    d_block_daemon_cp_element_group_236: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "d_block_daemon_cp_element_group_236"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= d_block_daemon_CP_6409_elements(234) & d_block_daemon_CP_6409_elements(235);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => d_block_daemon_CP_6409_elements(236), clk => clk, reset => reset); --
    end block;
    -- CP-element group 237:  transition  bypass 
    -- CP-element group 237: predecessors 
    -- CP-element group 237: 	8 
    -- CP-element group 237: successors 
    -- CP-element group 237:  members (1) 
      -- CP-element group 237: 	 branch_block_stmt_12832/merge_stmt_12918_dead_link/$entry
      -- 
    d_block_daemon_CP_6409_elements(237) <= d_block_daemon_CP_6409_elements(8);
    -- CP-element group 238:  fork  transition  output  bypass 
    -- CP-element group 238: predecessors 
    -- CP-element group 238: 	8 
    -- CP-element group 238: successors 
    -- CP-element group 238: 	239 
    -- CP-element group 238: 	240 
    -- CP-element group 238:  members (8) 
      -- CP-element group 238: 	 branch_block_stmt_12832/merge_stmt_12918__entry___PhiReq/phi_stmt_12919/phi_stmt_12919_sources/Interlock/Update/req
      -- CP-element group 238: 	 branch_block_stmt_12832/merge_stmt_12918__entry___PhiReq/phi_stmt_12919/phi_stmt_12919_sources/Interlock/Update/$entry
      -- CP-element group 238: 	 branch_block_stmt_12832/merge_stmt_12918__entry___PhiReq/phi_stmt_12919/phi_stmt_12919_sources/Interlock/Sample/req
      -- CP-element group 238: 	 branch_block_stmt_12832/merge_stmt_12918__entry___PhiReq/$entry
      -- CP-element group 238: 	 branch_block_stmt_12832/merge_stmt_12918__entry___PhiReq/phi_stmt_12919/phi_stmt_12919_sources/Interlock/Sample/$entry
      -- CP-element group 238: 	 branch_block_stmt_12832/merge_stmt_12918__entry___PhiReq/phi_stmt_12919/phi_stmt_12919_sources/Interlock/$entry
      -- CP-element group 238: 	 branch_block_stmt_12832/merge_stmt_12918__entry___PhiReq/phi_stmt_12919/phi_stmt_12919_sources/$entry
      -- CP-element group 238: 	 branch_block_stmt_12832/merge_stmt_12918__entry___PhiReq/phi_stmt_12919/$entry
      -- 
    req_7635_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7635_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_6409_elements(238), ack => countA_12863_12921_buf_req_0); -- 
    req_7640_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7640_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_6409_elements(238), ack => countA_12863_12921_buf_req_1); -- 
    d_block_daemon_CP_6409_elements(238) <= d_block_daemon_CP_6409_elements(8);
    -- CP-element group 239:  transition  input  bypass 
    -- CP-element group 239: predecessors 
    -- CP-element group 239: 	238 
    -- CP-element group 239: successors 
    -- CP-element group 239: 	241 
    -- CP-element group 239:  members (2) 
      -- CP-element group 239: 	 branch_block_stmt_12832/merge_stmt_12918__entry___PhiReq/phi_stmt_12919/phi_stmt_12919_sources/Interlock/Sample/ack
      -- CP-element group 239: 	 branch_block_stmt_12832/merge_stmt_12918__entry___PhiReq/phi_stmt_12919/phi_stmt_12919_sources/Interlock/Sample/$exit
      -- 
    ack_7636_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 239_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => countA_12863_12921_buf_ack_0, ack => d_block_daemon_CP_6409_elements(239)); -- 
    -- CP-element group 240:  transition  input  bypass 
    -- CP-element group 240: predecessors 
    -- CP-element group 240: 	238 
    -- CP-element group 240: successors 
    -- CP-element group 240: 	241 
    -- CP-element group 240:  members (2) 
      -- CP-element group 240: 	 branch_block_stmt_12832/merge_stmt_12918__entry___PhiReq/phi_stmt_12919/phi_stmt_12919_sources/Interlock/Update/ack
      -- CP-element group 240: 	 branch_block_stmt_12832/merge_stmt_12918__entry___PhiReq/phi_stmt_12919/phi_stmt_12919_sources/Interlock/Update/$exit
      -- 
    ack_7641_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 240_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => countA_12863_12921_buf_ack_1, ack => d_block_daemon_CP_6409_elements(240)); -- 
    -- CP-element group 241:  join  transition  output  bypass 
    -- CP-element group 241: predecessors 
    -- CP-element group 241: 	239 
    -- CP-element group 241: 	240 
    -- CP-element group 241: successors 
    -- CP-element group 241: 	246 
    -- CP-element group 241:  members (5) 
      -- CP-element group 241: 	 branch_block_stmt_12832/merge_stmt_12918__entry___PhiReq/phi_stmt_12919/phi_stmt_12919_req
      -- CP-element group 241: 	 branch_block_stmt_12832/merge_stmt_12918__entry___PhiReq/$exit
      -- CP-element group 241: 	 branch_block_stmt_12832/merge_stmt_12918__entry___PhiReq/phi_stmt_12919/phi_stmt_12919_sources/Interlock/$exit
      -- CP-element group 241: 	 branch_block_stmt_12832/merge_stmt_12918__entry___PhiReq/phi_stmt_12919/phi_stmt_12919_sources/$exit
      -- CP-element group 241: 	 branch_block_stmt_12832/merge_stmt_12918__entry___PhiReq/phi_stmt_12919/$exit
      -- 
    phi_stmt_12919_req_7642_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_12919_req_7642_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_6409_elements(241), ack => phi_stmt_12919_req_0); -- 
    d_block_daemon_cp_element_group_241: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "d_block_daemon_cp_element_group_241"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= d_block_daemon_CP_6409_elements(239) & d_block_daemon_CP_6409_elements(240);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => d_block_daemon_CP_6409_elements(241), clk => clk, reset => reset); --
    end block;
    -- CP-element group 242:  fork  transition  output  bypass 
    -- CP-element group 242: predecessors 
    -- CP-element group 242: 	209 
    -- CP-element group 242: successors 
    -- CP-element group 242: 	243 
    -- CP-element group 242: 	244 
    -- CP-element group 242:  members (8) 
      -- CP-element group 242: 	 branch_block_stmt_12832/NotGotNewKey_PhiReq/$entry
      -- CP-element group 242: 	 branch_block_stmt_12832/NotGotNewKey_PhiReq/phi_stmt_12919/phi_stmt_12919_sources/Interlock/Update/$entry
      -- CP-element group 242: 	 branch_block_stmt_12832/NotGotNewKey_PhiReq/phi_stmt_12919/phi_stmt_12919_sources/Interlock/Sample/req
      -- CP-element group 242: 	 branch_block_stmt_12832/NotGotNewKey_PhiReq/phi_stmt_12919/phi_stmt_12919_sources/Interlock/Update/req
      -- CP-element group 242: 	 branch_block_stmt_12832/NotGotNewKey_PhiReq/phi_stmt_12919/phi_stmt_12919_sources/Interlock/Sample/$entry
      -- CP-element group 242: 	 branch_block_stmt_12832/NotGotNewKey_PhiReq/phi_stmt_12919/phi_stmt_12919_sources/Interlock/$entry
      -- CP-element group 242: 	 branch_block_stmt_12832/NotGotNewKey_PhiReq/phi_stmt_12919/phi_stmt_12919_sources/$entry
      -- CP-element group 242: 	 branch_block_stmt_12832/NotGotNewKey_PhiReq/phi_stmt_12919/$entry
      -- 
    req_7658_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7658_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_6409_elements(242), ack => d_new_count_13047_12922_buf_req_0); -- 
    req_7663_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7663_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_6409_elements(242), ack => d_new_count_13047_12922_buf_req_1); -- 
    d_block_daemon_CP_6409_elements(242) <= d_block_daemon_CP_6409_elements(209);
    -- CP-element group 243:  transition  input  bypass 
    -- CP-element group 243: predecessors 
    -- CP-element group 243: 	242 
    -- CP-element group 243: successors 
    -- CP-element group 243: 	245 
    -- CP-element group 243:  members (2) 
      -- CP-element group 243: 	 branch_block_stmt_12832/NotGotNewKey_PhiReq/phi_stmt_12919/phi_stmt_12919_sources/Interlock/Sample/ack
      -- CP-element group 243: 	 branch_block_stmt_12832/NotGotNewKey_PhiReq/phi_stmt_12919/phi_stmt_12919_sources/Interlock/Sample/$exit
      -- 
    ack_7659_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 243_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_new_count_13047_12922_buf_ack_0, ack => d_block_daemon_CP_6409_elements(243)); -- 
    -- CP-element group 244:  transition  input  bypass 
    -- CP-element group 244: predecessors 
    -- CP-element group 244: 	242 
    -- CP-element group 244: successors 
    -- CP-element group 244: 	245 
    -- CP-element group 244:  members (2) 
      -- CP-element group 244: 	 branch_block_stmt_12832/NotGotNewKey_PhiReq/phi_stmt_12919/phi_stmt_12919_sources/Interlock/Update/$exit
      -- CP-element group 244: 	 branch_block_stmt_12832/NotGotNewKey_PhiReq/phi_stmt_12919/phi_stmt_12919_sources/Interlock/Update/ack
      -- 
    ack_7664_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 244_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_new_count_13047_12922_buf_ack_1, ack => d_block_daemon_CP_6409_elements(244)); -- 
    -- CP-element group 245:  join  transition  output  bypass 
    -- CP-element group 245: predecessors 
    -- CP-element group 245: 	243 
    -- CP-element group 245: 	244 
    -- CP-element group 245: successors 
    -- CP-element group 245: 	246 
    -- CP-element group 245:  members (5) 
      -- CP-element group 245: 	 branch_block_stmt_12832/NotGotNewKey_PhiReq/$exit
      -- CP-element group 245: 	 branch_block_stmt_12832/NotGotNewKey_PhiReq/phi_stmt_12919/phi_stmt_12919_sources/Interlock/$exit
      -- CP-element group 245: 	 branch_block_stmt_12832/NotGotNewKey_PhiReq/phi_stmt_12919/phi_stmt_12919_sources/$exit
      -- CP-element group 245: 	 branch_block_stmt_12832/NotGotNewKey_PhiReq/phi_stmt_12919/phi_stmt_12919_req
      -- CP-element group 245: 	 branch_block_stmt_12832/NotGotNewKey_PhiReq/phi_stmt_12919/$exit
      -- 
    phi_stmt_12919_req_7665_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_12919_req_7665_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => d_block_daemon_CP_6409_elements(245), ack => phi_stmt_12919_req_1); -- 
    d_block_daemon_cp_element_group_245: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "d_block_daemon_cp_element_group_245"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= d_block_daemon_CP_6409_elements(243) & d_block_daemon_CP_6409_elements(244);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => d_block_daemon_CP_6409_elements(245), clk => clk, reset => reset); --
    end block;
    -- CP-element group 246:  merge  place  bypass 
    -- CP-element group 246: predecessors 
    -- CP-element group 246: 	241 
    -- CP-element group 246: 	245 
    -- CP-element group 246: successors 
    -- CP-element group 246: 	247 
    -- CP-element group 246:  members (1) 
      -- CP-element group 246: 	 branch_block_stmt_12832/merge_stmt_12918_PhiReqMerge
      -- 
    d_block_daemon_CP_6409_elements(246) <= OrReduce(d_block_daemon_CP_6409_elements(241) & d_block_daemon_CP_6409_elements(245));
    -- CP-element group 247:  transition  bypass 
    -- CP-element group 247: predecessors 
    -- CP-element group 247: 	246 
    -- CP-element group 247: successors 
    -- CP-element group 247: 	248 
    -- CP-element group 247:  members (1) 
      -- CP-element group 247: 	 branch_block_stmt_12832/merge_stmt_12918_PhiAck/$entry
      -- 
    d_block_daemon_CP_6409_elements(247) <= d_block_daemon_CP_6409_elements(246);
    -- CP-element group 248:  transition  input  bypass 
    -- CP-element group 248: predecessors 
    -- CP-element group 248: 	247 
    -- CP-element group 248: successors 
    -- CP-element group 248: 	9 
    -- CP-element group 248:  members (2) 
      -- CP-element group 248: 	 branch_block_stmt_12832/merge_stmt_12918_PhiAck/$exit
      -- CP-element group 248: 	 branch_block_stmt_12832/merge_stmt_12918_PhiAck/phi_stmt_12919_ack
      -- 
    phi_stmt_12919_ack_7670_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 248_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_12919_ack_0, ack => d_block_daemon_CP_6409_elements(248)); -- 
    -- CP-element group 249:  join  transition  bypass  pipeline-parent 
    -- CP-element group 249: predecessors 
    -- CP-element group 249: 	71 
    -- CP-element group 249: 	183 
    -- CP-element group 249: successors 
    -- CP-element group 249: 	55 
    -- CP-element group 249:  members (2) 
      -- CP-element group 249: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/$exit
      -- CP-element group 249: 	 branch_block_stmt_12832/do_while_stmt_12924/do_while_stmt_12924_loop_body/phi_stmt_12926_phi_mux_ack_ps
      -- 
    d_block_daemon_cp_element_group_249: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 2,1 => 2);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "d_block_daemon_cp_element_group_249"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= d_block_daemon_CP_6409_elements(71) & d_block_daemon_CP_6409_elements(183);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => d_block_daemon_CP_6409_elements(249), clk => clk, reset => reset); --
    end block;
    do_while_stmt_12924_terminator_7375: loop_terminator -- 
      generic map (name => " do_while_stmt_12924_terminator_7375", max_iterations_in_flight =>2) 
      port map(loop_body_exit => d_block_daemon_CP_6409_elements(55),loop_continue => d_block_daemon_CP_6409_elements(192),loop_terminate => d_block_daemon_CP_6409_elements(190),loop_back => d_block_daemon_CP_6409_elements(53),loop_exit => d_block_daemon_CP_6409_elements(52),clk => clk, reset => reset); -- 
    phi_stmt_12926_phi_seq_6854_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= d_block_daemon_CP_6409_elements(66);
      d_block_daemon_CP_6409_elements(72)<= src_sample_reqs(0);
      src_sample_acks(0)  <= d_block_daemon_CP_6409_elements(72);
      d_block_daemon_CP_6409_elements(73)<= src_update_reqs(0);
      src_update_acks(0)  <= d_block_daemon_CP_6409_elements(74);
      d_block_daemon_CP_6409_elements(67) <= phi_mux_reqs(0);
      triggers(1)  <= d_block_daemon_CP_6409_elements(64);
      d_block_daemon_CP_6409_elements(76)<= src_sample_reqs(1);
      src_sample_acks(1)  <= d_block_daemon_CP_6409_elements(78);
      d_block_daemon_CP_6409_elements(77)<= src_update_reqs(1);
      src_update_acks(1)  <= d_block_daemon_CP_6409_elements(79);
      d_block_daemon_CP_6409_elements(65) <= phi_mux_reqs(1);
      phi_stmt_12926_phi_seq_6854 : phi_sequencer_v2-- 
        generic map (place_capacity => 2, ntriggers => 2, name => "phi_stmt_12926_phi_seq_6854") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => d_block_daemon_CP_6409_elements(60), 
          phi_sample_ack => d_block_daemon_CP_6409_elements(62), 
          phi_update_req => d_block_daemon_CP_6409_elements(61), 
          phi_update_ack => d_block_daemon_CP_6409_elements(63), 
          phi_mux_ack => d_block_daemon_CP_6409_elements(71), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_6805_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= d_block_daemon_CP_6409_elements(56);
        preds(1)  <= d_block_daemon_CP_6409_elements(57);
        entry_tmerge_6805 : transition_merge -- 
          generic map(name => " entry_tmerge_6805")
          port map (preds => preds, symbol_out => d_block_daemon_CP_6409_elements(58));
          -- 
    end block;
    phi_stmt_12926_req_merge_6825_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= d_block_daemon_CP_6409_elements(69);
        preds(1)  <= d_block_daemon_CP_6409_elements(70);
        phi_stmt_12926_req_merge_6825 : transition_merge -- 
          generic map(name => " phi_stmt_12926_req_merge_6825")
          port map (preds => preds, symbol_out => d_block_daemon_CP_6409_elements(68));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal EQ_u1_u1_12855_wire : std_logic_vector(0 downto 0);
    signal EQ_u1_u1_13055_wire : std_logic_vector(0 downto 0);
    signal K0_12859 : std_logic_vector(127 downto 0);
    signal K0_12985_delayed_10_13016 : std_logic_vector(127 downto 0);
    signal K10_12917 : std_logic_vector(127 downto 0);
    signal K10_12936_delayed_1_12936 : std_logic_vector(127 downto 0);
    signal K1_12872 : std_logic_vector(127 downto 0);
    signal K1_12980_delayed_9_13008 : std_logic_vector(127 downto 0);
    signal K2_12877 : std_logic_vector(127 downto 0);
    signal K2_12975_delayed_8_13000 : std_logic_vector(127 downto 0);
    signal K3_12882 : std_logic_vector(127 downto 0);
    signal K3_12970_delayed_7_12992 : std_logic_vector(127 downto 0);
    signal K4_12887 : std_logic_vector(127 downto 0);
    signal K4_12965_delayed_6_12984 : std_logic_vector(127 downto 0);
    signal K5_12892 : std_logic_vector(127 downto 0);
    signal K5_12960_delayed_5_12976 : std_logic_vector(127 downto 0);
    signal K6_12897 : std_logic_vector(127 downto 0);
    signal K6_12955_delayed_4_12968 : std_logic_vector(127 downto 0);
    signal K7_12902 : std_logic_vector(127 downto 0);
    signal K7_12950_delayed_3_12960 : std_logic_vector(127 downto 0);
    signal K8_12907 : std_logic_vector(127 downto 0);
    signal K8_12945_delayed_2_12952 : std_logic_vector(127 downto 0);
    signal K9_12912 : std_logic_vector(127 downto 0);
    signal K9_12940_delayed_1_12944 : std_logic_vector(127 downto 0);
    signal RConstant_10_12912 : std_logic_vector(7 downto 0);
    signal RConstant_11_12917 : std_logic_vector(7 downto 0);
    signal RConstant_2_12872 : std_logic_vector(7 downto 0);
    signal RConstant_3_12877 : std_logic_vector(7 downto 0);
    signal RConstant_4_12882 : std_logic_vector(7 downto 0);
    signal RConstant_5_12887 : std_logic_vector(7 downto 0);
    signal RConstant_6_12892 : std_logic_vector(7 downto 0);
    signal RConstant_7_12897 : std_logic_vector(7 downto 0);
    signal RConstant_8_12902 : std_logic_vector(7 downto 0);
    signal RConstant_9_12907 : std_logic_vector(7 downto 0);
    signal R_LAST_12947_wire_constant : std_logic_vector(0 downto 0);
    signal R_NOT_LAST_12955_wire_constant : std_logic_vector(0 downto 0);
    signal R_NOT_LAST_12963_wire_constant : std_logic_vector(0 downto 0);
    signal R_NOT_LAST_12971_wire_constant : std_logic_vector(0 downto 0);
    signal R_NOT_LAST_12979_wire_constant : std_logic_vector(0 downto 0);
    signal R_NOT_LAST_12987_wire_constant : std_logic_vector(0 downto 0);
    signal R_NOT_LAST_12995_wire_constant : std_logic_vector(0 downto 0);
    signal R_NOT_LAST_13003_wire_constant : std_logic_vector(0 downto 0);
    signal R_NOT_LAST_13011_wire_constant : std_logic_vector(0 downto 0);
    signal R_NOT_LAST_13019_wire_constant : std_logic_vector(0 downto 0);
    signal R_RConstant_1_12869_wire_constant : std_logic_vector(7 downto 0);
    signal R_ZERO_COUNT_12928_wire_constant : std_logic_vector(14 downto 0);
    signal ULT_u15_u1_13033_wire : std_logic_vector(0 downto 0);
    signal countA_12863 : std_logic_vector(14 downto 0);
    signal countA_12863_12921_buffered : std_logic_vector(14 downto 0);
    signal countB_12919 : std_logic_vector(14 downto 0);
    signal count_var_12926 : std_logic_vector(14 downto 0);
    signal d_get_key_12843 : std_logic_vector(0 downto 0);
    signal d_get_new_key_13043 : std_logic_vector(0 downto 0);
    signal d_init_cmd_12839 : std_logic_vector(143 downto 0);
    signal d_init_count_12847 : std_logic_vector(14 downto 0);
    signal d_init_count_12847_12865_buffered : std_logic_vector(14 downto 0);
    signal d_init_key_12851 : std_logic_vector(127 downto 0);
    signal d_init_key_12851_12861_buffered : std_logic_vector(127 downto 0);
    signal d_new_cmd_13039 : std_logic_vector(143 downto 0);
    signal d_new_count_13047 : std_logic_vector(14 downto 0);
    signal d_new_count_13047_12866_buffered : std_logic_vector(14 downto 0);
    signal d_new_count_13047_12922_buffered : std_logic_vector(14 downto 0);
    signal d_new_key_13051 : std_logic_vector(127 downto 0);
    signal d_new_key_13051_12862_buffered : std_logic_vector(127 downto 0);
    signal in128_12933 : std_logic_vector(127 downto 0);
    signal konst_12834_wire_constant : std_logic_vector(0 downto 0);
    signal konst_12854_wire_constant : std_logic_vector(0 downto 0);
    signal konst_13027_wire_constant : std_logic_vector(14 downto 0);
    signal konst_13035_wire_constant : std_logic_vector(0 downto 0);
    signal konst_13054_wire_constant : std_logic_vector(0 downto 0);
    signal n_count_var_13029 : std_logic_vector(14 downto 0);
    signal n_count_var_13029_12929_buffered : std_logic_vector(14 downto 0);
    signal round_S0_13021 : std_logic_vector(127 downto 0);
    signal round_S10_12941 : std_logic_vector(127 downto 0);
    signal round_S1_13013 : std_logic_vector(127 downto 0);
    signal round_S2_13005 : std_logic_vector(127 downto 0);
    signal round_S3_12997 : std_logic_vector(127 downto 0);
    signal round_S4_12989 : std_logic_vector(127 downto 0);
    signal round_S5_12981 : std_logic_vector(127 downto 0);
    signal round_S6_12973 : std_logic_vector(127 downto 0);
    signal round_S7_12965 : std_logic_vector(127 downto 0);
    signal round_S8_12957 : std_logic_vector(127 downto 0);
    signal round_S9_12949 : std_logic_vector(127 downto 0);
    signal xxd_block_daemonxxLAST : std_logic_vector(0 downto 0);
    signal xxd_block_daemonxxNOT_LAST : std_logic_vector(0 downto 0);
    signal xxd_block_daemonxxRConstant_1 : std_logic_vector(7 downto 0);
    signal xxd_block_daemonxxZERO_COUNT : std_logic_vector(14 downto 0);
    -- 
  begin -- 
    R_LAST_12947_wire_constant <= "1";
    R_NOT_LAST_12955_wire_constant <= "0";
    R_NOT_LAST_12963_wire_constant <= "0";
    R_NOT_LAST_12971_wire_constant <= "0";
    R_NOT_LAST_12979_wire_constant <= "0";
    R_NOT_LAST_12987_wire_constant <= "0";
    R_NOT_LAST_12995_wire_constant <= "0";
    R_NOT_LAST_13003_wire_constant <= "0";
    R_NOT_LAST_13011_wire_constant <= "0";
    R_NOT_LAST_13019_wire_constant <= "0";
    R_RConstant_1_12869_wire_constant <= "00000001";
    R_ZERO_COUNT_12928_wire_constant <= "000000000000000";
    konst_12834_wire_constant <= "1";
    konst_12854_wire_constant <= "0";
    konst_13027_wire_constant <= "000000000000001";
    konst_13035_wire_constant <= "1";
    konst_13054_wire_constant <= "1";
    xxd_block_daemonxxLAST <= "1";
    xxd_block_daemonxxNOT_LAST <= "0";
    xxd_block_daemonxxRConstant_1 <= "00000001";
    xxd_block_daemonxxZERO_COUNT <= "000000000000000";
    phi_stmt_12859: Block -- phi operator 
      signal idata: std_logic_vector(255 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= d_init_key_12851_12861_buffered & d_new_key_13051_12862_buffered;
      req <= phi_stmt_12859_req_0 & phi_stmt_12859_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_12859",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 128) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_12859_ack_0,
          idata => idata,
          odata => K0_12859,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_12859
    phi_stmt_12863: Block -- phi operator 
      signal idata: std_logic_vector(29 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= d_init_count_12847_12865_buffered & d_new_count_13047_12866_buffered;
      req <= phi_stmt_12863_req_0 & phi_stmt_12863_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_12863",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 15) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_12863_ack_0,
          idata => idata,
          odata => countA_12863,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_12863
    phi_stmt_12919: Block -- phi operator 
      signal idata: std_logic_vector(29 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= countA_12863_12921_buffered & d_new_count_13047_12922_buffered;
      req <= phi_stmt_12919_req_0 & phi_stmt_12919_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_12919",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 15) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_12919_ack_0,
          idata => idata,
          odata => countB_12919,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_12919
    phi_stmt_12926: Block -- phi operator 
      signal idata: std_logic_vector(29 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_COUNT_12928_wire_constant & n_count_var_13029_12929_buffered;
      req <= phi_stmt_12926_req_0 & phi_stmt_12926_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_12926",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 15) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_12926_ack_0,
          idata => idata,
          odata => count_var_12926,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_12926
    -- flow-through slice operator slice_12842_inst
    d_get_key_12843 <= d_init_cmd_12839(143 downto 143);
    -- flow-through slice operator slice_12846_inst
    d_init_count_12847 <= d_init_cmd_12839(142 downto 128);
    -- flow-through slice operator slice_12850_inst
    d_init_key_12851 <= d_init_cmd_12839(127 downto 0);
    -- flow-through slice operator slice_13042_inst
    d_get_new_key_13043 <= d_new_cmd_13039(143 downto 143);
    -- flow-through slice operator slice_13046_inst
    d_new_count_13047 <= d_new_cmd_13039(142 downto 128);
    -- flow-through slice operator slice_13050_inst
    d_new_key_13051 <= d_new_cmd_13039(127 downto 0);
    W_K0_12985_delayed_10_13014_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_K0_12985_delayed_10_13014_inst_req_0;
      W_K0_12985_delayed_10_13014_inst_ack_0<= wack(0);
      rreq(0) <= W_K0_12985_delayed_10_13014_inst_req_1;
      W_K0_12985_delayed_10_13014_inst_ack_1<= rack(0);
      W_K0_12985_delayed_10_13014_inst : InterlockBuffer generic map ( -- 
        name => "W_K0_12985_delayed_10_13014_inst",
        buffer_size => 10,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 128,
        out_data_width => 128,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => K0_12859,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => K0_12985_delayed_10_13016,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_K10_12936_delayed_1_12934_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_K10_12936_delayed_1_12934_inst_req_0;
      W_K10_12936_delayed_1_12934_inst_ack_0<= wack(0);
      rreq(0) <= W_K10_12936_delayed_1_12934_inst_req_1;
      W_K10_12936_delayed_1_12934_inst_ack_1<= rack(0);
      W_K10_12936_delayed_1_12934_inst : InterlockBuffer generic map ( -- 
        name => "W_K10_12936_delayed_1_12934_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 128,
        out_data_width => 128,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => K10_12917,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => K10_12936_delayed_1_12936,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_K1_12980_delayed_9_13006_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_K1_12980_delayed_9_13006_inst_req_0;
      W_K1_12980_delayed_9_13006_inst_ack_0<= wack(0);
      rreq(0) <= W_K1_12980_delayed_9_13006_inst_req_1;
      W_K1_12980_delayed_9_13006_inst_ack_1<= rack(0);
      W_K1_12980_delayed_9_13006_inst : InterlockBuffer generic map ( -- 
        name => "W_K1_12980_delayed_9_13006_inst",
        buffer_size => 9,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 128,
        out_data_width => 128,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => K1_12872,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => K1_12980_delayed_9_13008,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_K2_12975_delayed_8_12998_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_K2_12975_delayed_8_12998_inst_req_0;
      W_K2_12975_delayed_8_12998_inst_ack_0<= wack(0);
      rreq(0) <= W_K2_12975_delayed_8_12998_inst_req_1;
      W_K2_12975_delayed_8_12998_inst_ack_1<= rack(0);
      W_K2_12975_delayed_8_12998_inst : InterlockBuffer generic map ( -- 
        name => "W_K2_12975_delayed_8_12998_inst",
        buffer_size => 8,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 128,
        out_data_width => 128,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => K2_12877,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => K2_12975_delayed_8_13000,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_K3_12970_delayed_7_12990_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_K3_12970_delayed_7_12990_inst_req_0;
      W_K3_12970_delayed_7_12990_inst_ack_0<= wack(0);
      rreq(0) <= W_K3_12970_delayed_7_12990_inst_req_1;
      W_K3_12970_delayed_7_12990_inst_ack_1<= rack(0);
      W_K3_12970_delayed_7_12990_inst : InterlockBuffer generic map ( -- 
        name => "W_K3_12970_delayed_7_12990_inst",
        buffer_size => 7,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 128,
        out_data_width => 128,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => K3_12882,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => K3_12970_delayed_7_12992,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_K4_12965_delayed_6_12982_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_K4_12965_delayed_6_12982_inst_req_0;
      W_K4_12965_delayed_6_12982_inst_ack_0<= wack(0);
      rreq(0) <= W_K4_12965_delayed_6_12982_inst_req_1;
      W_K4_12965_delayed_6_12982_inst_ack_1<= rack(0);
      W_K4_12965_delayed_6_12982_inst : InterlockBuffer generic map ( -- 
        name => "W_K4_12965_delayed_6_12982_inst",
        buffer_size => 6,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 128,
        out_data_width => 128,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => K4_12887,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => K4_12965_delayed_6_12984,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_K5_12960_delayed_5_12974_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_K5_12960_delayed_5_12974_inst_req_0;
      W_K5_12960_delayed_5_12974_inst_ack_0<= wack(0);
      rreq(0) <= W_K5_12960_delayed_5_12974_inst_req_1;
      W_K5_12960_delayed_5_12974_inst_ack_1<= rack(0);
      W_K5_12960_delayed_5_12974_inst : InterlockBuffer generic map ( -- 
        name => "W_K5_12960_delayed_5_12974_inst",
        buffer_size => 5,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 128,
        out_data_width => 128,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => K5_12892,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => K5_12960_delayed_5_12976,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_K6_12955_delayed_4_12966_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_K6_12955_delayed_4_12966_inst_req_0;
      W_K6_12955_delayed_4_12966_inst_ack_0<= wack(0);
      rreq(0) <= W_K6_12955_delayed_4_12966_inst_req_1;
      W_K6_12955_delayed_4_12966_inst_ack_1<= rack(0);
      W_K6_12955_delayed_4_12966_inst : InterlockBuffer generic map ( -- 
        name => "W_K6_12955_delayed_4_12966_inst",
        buffer_size => 4,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 128,
        out_data_width => 128,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => K6_12897,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => K6_12955_delayed_4_12968,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_K7_12950_delayed_3_12958_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_K7_12950_delayed_3_12958_inst_req_0;
      W_K7_12950_delayed_3_12958_inst_ack_0<= wack(0);
      rreq(0) <= W_K7_12950_delayed_3_12958_inst_req_1;
      W_K7_12950_delayed_3_12958_inst_ack_1<= rack(0);
      W_K7_12950_delayed_3_12958_inst : InterlockBuffer generic map ( -- 
        name => "W_K7_12950_delayed_3_12958_inst",
        buffer_size => 3,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 128,
        out_data_width => 128,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => K7_12902,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => K7_12950_delayed_3_12960,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_K8_12945_delayed_2_12950_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_K8_12945_delayed_2_12950_inst_req_0;
      W_K8_12945_delayed_2_12950_inst_ack_0<= wack(0);
      rreq(0) <= W_K8_12945_delayed_2_12950_inst_req_1;
      W_K8_12945_delayed_2_12950_inst_ack_1<= rack(0);
      W_K8_12945_delayed_2_12950_inst : InterlockBuffer generic map ( -- 
        name => "W_K8_12945_delayed_2_12950_inst",
        buffer_size => 2,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 128,
        out_data_width => 128,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => K8_12907,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => K8_12945_delayed_2_12952,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_K9_12940_delayed_1_12942_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_K9_12940_delayed_1_12942_inst_req_0;
      W_K9_12940_delayed_1_12942_inst_ack_0<= wack(0);
      rreq(0) <= W_K9_12940_delayed_1_12942_inst_req_1;
      W_K9_12940_delayed_1_12942_inst_ack_1<= rack(0);
      W_K9_12940_delayed_1_12942_inst : InterlockBuffer generic map ( -- 
        name => "W_K9_12940_delayed_1_12942_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 128,
        out_data_width => 128,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => K9_12912,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => K9_12940_delayed_1_12944,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    countA_12863_12921_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= countA_12863_12921_buf_req_0;
      countA_12863_12921_buf_ack_0<= wack(0);
      rreq(0) <= countA_12863_12921_buf_req_1;
      countA_12863_12921_buf_ack_1<= rack(0);
      countA_12863_12921_buf : InterlockBuffer generic map ( -- 
        name => "countA_12863_12921_buf",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 15,
        out_data_width => 15,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => countA_12863,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => countA_12863_12921_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    d_init_count_12847_12865_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= d_init_count_12847_12865_buf_req_0;
      d_init_count_12847_12865_buf_ack_0<= wack(0);
      rreq(0) <= d_init_count_12847_12865_buf_req_1;
      d_init_count_12847_12865_buf_ack_1<= rack(0);
      d_init_count_12847_12865_buf : InterlockBuffer generic map ( -- 
        name => "d_init_count_12847_12865_buf",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 15,
        out_data_width => 15,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => d_init_count_12847,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => d_init_count_12847_12865_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    d_init_key_12851_12861_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= d_init_key_12851_12861_buf_req_0;
      d_init_key_12851_12861_buf_ack_0<= wack(0);
      rreq(0) <= d_init_key_12851_12861_buf_req_1;
      d_init_key_12851_12861_buf_ack_1<= rack(0);
      d_init_key_12851_12861_buf : InterlockBuffer generic map ( -- 
        name => "d_init_key_12851_12861_buf",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 128,
        out_data_width => 128,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => d_init_key_12851,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => d_init_key_12851_12861_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    d_new_count_13047_12866_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= d_new_count_13047_12866_buf_req_0;
      d_new_count_13047_12866_buf_ack_0<= wack(0);
      rreq(0) <= d_new_count_13047_12866_buf_req_1;
      d_new_count_13047_12866_buf_ack_1<= rack(0);
      d_new_count_13047_12866_buf : InterlockBuffer generic map ( -- 
        name => "d_new_count_13047_12866_buf",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 15,
        out_data_width => 15,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => d_new_count_13047,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => d_new_count_13047_12866_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    d_new_count_13047_12922_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= d_new_count_13047_12922_buf_req_0;
      d_new_count_13047_12922_buf_ack_0<= wack(0);
      rreq(0) <= d_new_count_13047_12922_buf_req_1;
      d_new_count_13047_12922_buf_ack_1<= rack(0);
      d_new_count_13047_12922_buf : InterlockBuffer generic map ( -- 
        name => "d_new_count_13047_12922_buf",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 15,
        out_data_width => 15,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => d_new_count_13047,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => d_new_count_13047_12922_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    d_new_key_13051_12862_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= d_new_key_13051_12862_buf_req_0;
      d_new_key_13051_12862_buf_ack_0<= wack(0);
      rreq(0) <= d_new_key_13051_12862_buf_req_1;
      d_new_key_13051_12862_buf_ack_1<= rack(0);
      d_new_key_13051_12862_buf : InterlockBuffer generic map ( -- 
        name => "d_new_key_13051_12862_buf",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 128,
        out_data_width => 128,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => d_new_key_13051,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => d_new_key_13051_12862_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_count_var_13029_12929_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_count_var_13029_12929_buf_req_0;
      n_count_var_13029_12929_buf_ack_0<= wack(0);
      rreq(0) <= n_count_var_13029_12929_buf_req_1;
      n_count_var_13029_12929_buf_ack_1<= rack(0);
      n_count_var_13029_12929_buf : InterlockBuffer generic map ( -- 
        name => "n_count_var_13029_12929_buf",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 15,
        out_data_width => 15,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_count_var_13029,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_count_var_13029_12929_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    do_while_stmt_12924_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= ULT_u15_u1_13033_wire;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_12924_branch", condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_12924_branch_req_0,
          ack0 => do_while_stmt_12924_branch_ack_0,
          ack1 => do_while_stmt_12924_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_12852_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= EQ_u1_u1_12855_wire;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_12852_branch", condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_12852_branch_req_0,
          ack0 => if_stmt_12852_branch_ack_0,
          ack1 => if_stmt_12852_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_13052_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= EQ_u1_u1_13055_wire;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_13052_branch", condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_13052_branch_req_0,
          ack0 => if_stmt_13052_branch_ack_0,
          ack1 => if_stmt_13052_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- shared split operator group (0) : ADD_u15_u15_13028_inst 
    ApIntAdd_group_0: Block -- 
      signal data_in: std_logic_vector(14 downto 0);
      signal data_out: std_logic_vector(14 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= count_var_12926;
      n_count_var_13029 <= data_out(14 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u15_u15_13028_inst_req_0;
      ADD_u15_u15_13028_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u15_u15_13028_inst_req_1;
      ADD_u15_u15_13028_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(name => "gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_0",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 15,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 15,
          constant_operand => "000000000000001",
          constant_width => 15,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- binary operator EQ_u1_u1_12855_inst
    process(d_get_key_12843) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(d_get_key_12843, konst_12854_wire_constant, tmp_var);
      EQ_u1_u1_12855_wire <= tmp_var; -- 
    end process;
    -- binary operator EQ_u1_u1_13055_inst
    process(d_get_new_key_13043) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(d_get_new_key_13043, konst_13054_wire_constant, tmp_var);
      EQ_u1_u1_13055_wire <= tmp_var; -- 
    end process;
    -- binary operator ULT_u15_u1_13033_inst
    process(n_count_var_13029, countB_12919) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(n_count_var_13029, countB_12919, tmp_var);
      ULT_u15_u1_13033_wire <= tmp_var; -- 
    end process;
    -- binary operator XOR_u128_u128_12940_inst
    process(in128_12933, K10_12936_delayed_1_12936) -- 
      variable tmp_var : std_logic_vector(127 downto 0); -- 
    begin -- 
      ApIntXor_proc(in128_12933, K10_12936_delayed_1_12936, tmp_var);
      round_S10_12941 <= tmp_var; -- 
    end process;
    -- shared inport operator group (0) : RPIPE_d_cmd_pipe_12838_inst RPIPE_d_cmd_pipe_13038_inst 
    InportGroup0: Block -- 
      signal data_out: std_logic_vector(287 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 1 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= RPIPE_d_cmd_pipe_12838_inst_req_0;
      reqL_unguarded(0) <= RPIPE_d_cmd_pipe_13038_inst_req_0;
      RPIPE_d_cmd_pipe_12838_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_d_cmd_pipe_13038_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= RPIPE_d_cmd_pipe_12838_inst_req_1;
      reqR_unguarded(0) <= RPIPE_d_cmd_pipe_13038_inst_req_1;
      RPIPE_d_cmd_pipe_12838_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_d_cmd_pipe_13038_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      gI: SplitGuardInterface generic map(name => "gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      d_init_cmd_12839 <= data_out(287 downto 144);
      d_new_cmd_13039 <= data_out(143 downto 0);
      d_cmd_pipe_read_0: InputPortRevised -- 
        generic map ( name => "d_cmd_pipe_read_0", data_width => 144,  num_reqs => 2,  output_buffering => outBUFs,   no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => d_cmd_pipe_pipe_read_req(0),
          oack => d_cmd_pipe_pipe_read_ack(0),
          odata => d_cmd_pipe_pipe_read_data(143 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared inport operator group (1) : RPIPE_d_in_buf_12932_inst 
    InportGroup1: Block -- 
      signal data_out: std_logic_vector(127 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_d_in_buf_12932_inst_req_0;
      RPIPE_d_in_buf_12932_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_d_in_buf_12932_inst_req_1;
      RPIPE_d_in_buf_12932_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      gI: SplitGuardInterface generic map(name => "gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      in128_12933 <= data_out(127 downto 0);
      d_in_buf_read_1: InputPortRevised -- 
        generic map ( name => "d_in_buf_read_1", data_width => 128,  num_reqs => 1,  output_buffering => outBUFs,   no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => d_in_buf_pipe_read_req(0),
          oack => d_in_buf_pipe_read_ack(0),
          odata => d_in_buf_pipe_read_data(127 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 1
    -- shared outport operator group (0) : WPIPE_d_block_done_12833_inst WPIPE_d_block_done_13034_inst 
    OutportGroup0: Block -- 
      signal data_in: std_logic_vector(1 downto 0);
      signal sample_req, sample_ack : BooleanArray( 1 downto 0);
      signal update_req, update_ack : BooleanArray( 1 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 1 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      sample_req_unguarded(1) <= WPIPE_d_block_done_12833_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_d_block_done_13034_inst_req_0;
      WPIPE_d_block_done_12833_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_d_block_done_13034_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(1) <= WPIPE_d_block_done_12833_inst_req_1;
      update_req_unguarded(0) <= WPIPE_d_block_done_13034_inst_req_1;
      WPIPE_d_block_done_12833_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_d_block_done_13034_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      gI: SplitGuardInterface generic map(name => "gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      data_in <= konst_12834_wire_constant & konst_13035_wire_constant;
      d_block_done_write_0: OutputPortRevised -- 
        generic map ( name => "d_block_done", data_width => 1, num_reqs => 2, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => d_block_done_pipe_write_req(0),
          oack => d_block_done_pipe_write_ack(0),
          odata => d_block_done_pipe_write_data(0 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_d_out_buf_13022_inst 
    OutportGroup1: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_d_out_buf_13022_inst_req_0;
      WPIPE_d_out_buf_13022_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_d_out_buf_13022_inst_req_1;
      WPIPE_d_out_buf_13022_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      gI: SplitGuardInterface generic map(name => "gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      data_in <= round_S0_13021;
      d_out_buf_write_1: OutputPortRevised -- 
        generic map ( name => "d_out_buf", data_width => 128, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => d_out_buf_pipe_write_req(0),
          oack => d_out_buf_pipe_write_ack(0),
          odata => d_out_buf_pipe_write_data(127 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared call operator group (0) : call_stmt_12917_call call_stmt_12912_call call_stmt_12907_call call_stmt_12902_call call_stmt_12897_call call_stmt_12892_call call_stmt_12887_call call_stmt_12882_call call_stmt_12877_call call_stmt_12872_call 
    key_expand_single_call_group_0: Block -- 
      signal data_in: std_logic_vector(1359 downto 0);
      signal data_out: std_logic_vector(1359 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 9 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 9 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 9 downto 0);
      signal guard_vector : std_logic_vector( 9 downto 0);
      constant inBUFs : IntegerArray(9 downto 0) := (9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(9 downto 0) := (9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(9 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false);
      constant guardBuffering: IntegerArray(9 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2);
      -- 
    begin -- 
      reqL_unguarded(9) <= call_stmt_12917_call_req_0;
      reqL_unguarded(8) <= call_stmt_12912_call_req_0;
      reqL_unguarded(7) <= call_stmt_12907_call_req_0;
      reqL_unguarded(6) <= call_stmt_12902_call_req_0;
      reqL_unguarded(5) <= call_stmt_12897_call_req_0;
      reqL_unguarded(4) <= call_stmt_12892_call_req_0;
      reqL_unguarded(3) <= call_stmt_12887_call_req_0;
      reqL_unguarded(2) <= call_stmt_12882_call_req_0;
      reqL_unguarded(1) <= call_stmt_12877_call_req_0;
      reqL_unguarded(0) <= call_stmt_12872_call_req_0;
      call_stmt_12917_call_ack_0 <= ackL_unguarded(9);
      call_stmt_12912_call_ack_0 <= ackL_unguarded(8);
      call_stmt_12907_call_ack_0 <= ackL_unguarded(7);
      call_stmt_12902_call_ack_0 <= ackL_unguarded(6);
      call_stmt_12897_call_ack_0 <= ackL_unguarded(5);
      call_stmt_12892_call_ack_0 <= ackL_unguarded(4);
      call_stmt_12887_call_ack_0 <= ackL_unguarded(3);
      call_stmt_12882_call_ack_0 <= ackL_unguarded(2);
      call_stmt_12877_call_ack_0 <= ackL_unguarded(1);
      call_stmt_12872_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(9) <= call_stmt_12917_call_req_1;
      reqR_unguarded(8) <= call_stmt_12912_call_req_1;
      reqR_unguarded(7) <= call_stmt_12907_call_req_1;
      reqR_unguarded(6) <= call_stmt_12902_call_req_1;
      reqR_unguarded(5) <= call_stmt_12897_call_req_1;
      reqR_unguarded(4) <= call_stmt_12892_call_req_1;
      reqR_unguarded(3) <= call_stmt_12887_call_req_1;
      reqR_unguarded(2) <= call_stmt_12882_call_req_1;
      reqR_unguarded(1) <= call_stmt_12877_call_req_1;
      reqR_unguarded(0) <= call_stmt_12872_call_req_1;
      call_stmt_12917_call_ack_1 <= ackR_unguarded(9);
      call_stmt_12912_call_ack_1 <= ackR_unguarded(8);
      call_stmt_12907_call_ack_1 <= ackR_unguarded(7);
      call_stmt_12902_call_ack_1 <= ackR_unguarded(6);
      call_stmt_12897_call_ack_1 <= ackR_unguarded(5);
      call_stmt_12892_call_ack_1 <= ackR_unguarded(4);
      call_stmt_12887_call_ack_1 <= ackR_unguarded(3);
      call_stmt_12882_call_ack_1 <= ackR_unguarded(2);
      call_stmt_12877_call_ack_1 <= ackR_unguarded(1);
      call_stmt_12872_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      key_expand_single_call_group_0_accessRegulator_0: access_regulator_base generic map (name => "key_expand_single_call_group_0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      key_expand_single_call_group_0_accessRegulator_1: access_regulator_base generic map (name => "key_expand_single_call_group_0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      key_expand_single_call_group_0_accessRegulator_2: access_regulator_base generic map (name => "key_expand_single_call_group_0_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      key_expand_single_call_group_0_accessRegulator_3: access_regulator_base generic map (name => "key_expand_single_call_group_0_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      key_expand_single_call_group_0_accessRegulator_4: access_regulator_base generic map (name => "key_expand_single_call_group_0_accessRegulator_4", num_slots => 1) -- 
        port map (req => reqL_unregulated(4), -- 
          ack => ackL_unregulated(4),
          regulated_req => reqL(4),
          regulated_ack => ackL(4),
          release_req => reqR(4),
          release_ack => ackR(4),
          clk => clk, reset => reset); -- 
      key_expand_single_call_group_0_accessRegulator_5: access_regulator_base generic map (name => "key_expand_single_call_group_0_accessRegulator_5", num_slots => 1) -- 
        port map (req => reqL_unregulated(5), -- 
          ack => ackL_unregulated(5),
          regulated_req => reqL(5),
          regulated_ack => ackL(5),
          release_req => reqR(5),
          release_ack => ackR(5),
          clk => clk, reset => reset); -- 
      key_expand_single_call_group_0_accessRegulator_6: access_regulator_base generic map (name => "key_expand_single_call_group_0_accessRegulator_6", num_slots => 1) -- 
        port map (req => reqL_unregulated(6), -- 
          ack => ackL_unregulated(6),
          regulated_req => reqL(6),
          regulated_ack => ackL(6),
          release_req => reqR(6),
          release_ack => ackR(6),
          clk => clk, reset => reset); -- 
      key_expand_single_call_group_0_accessRegulator_7: access_regulator_base generic map (name => "key_expand_single_call_group_0_accessRegulator_7", num_slots => 1) -- 
        port map (req => reqL_unregulated(7), -- 
          ack => ackL_unregulated(7),
          regulated_req => reqL(7),
          regulated_ack => ackL(7),
          release_req => reqR(7),
          release_ack => ackR(7),
          clk => clk, reset => reset); -- 
      key_expand_single_call_group_0_accessRegulator_8: access_regulator_base generic map (name => "key_expand_single_call_group_0_accessRegulator_8", num_slots => 1) -- 
        port map (req => reqL_unregulated(8), -- 
          ack => ackL_unregulated(8),
          regulated_req => reqL(8),
          regulated_ack => ackL(8),
          release_req => reqR(8),
          release_ack => ackR(8),
          clk => clk, reset => reset); -- 
      key_expand_single_call_group_0_accessRegulator_9: access_regulator_base generic map (name => "key_expand_single_call_group_0_accessRegulator_9", num_slots => 1) -- 
        port map (req => reqL_unregulated(9), -- 
          ack => ackL_unregulated(9),
          regulated_req => reqL(9),
          regulated_ack => ackL(9),
          release_req => reqR(9),
          release_ack => ackR(9),
          clk => clk, reset => reset); -- 
      gI: SplitGuardInterface generic map(name => "gI", nreqs => 10, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= K9_12912 & RConstant_10_12912 & K8_12907 & RConstant_9_12907 & K7_12902 & RConstant_8_12902 & K6_12897 & RConstant_7_12897 & K5_12892 & RConstant_6_12892 & K4_12887 & RConstant_5_12887 & K3_12882 & RConstant_4_12882 & K2_12877 & RConstant_3_12877 & K1_12872 & RConstant_2_12872 & K0_12859 & R_RConstant_1_12869_wire_constant;
      K10_12917 <= data_out(1359 downto 1232);
      RConstant_11_12917 <= data_out(1231 downto 1224);
      K9_12912 <= data_out(1223 downto 1096);
      RConstant_10_12912 <= data_out(1095 downto 1088);
      K8_12907 <= data_out(1087 downto 960);
      RConstant_9_12907 <= data_out(959 downto 952);
      K7_12902 <= data_out(951 downto 824);
      RConstant_8_12902 <= data_out(823 downto 816);
      K6_12897 <= data_out(815 downto 688);
      RConstant_7_12897 <= data_out(687 downto 680);
      K5_12892 <= data_out(679 downto 552);
      RConstant_6_12892 <= data_out(551 downto 544);
      K4_12887 <= data_out(543 downto 416);
      RConstant_5_12887 <= data_out(415 downto 408);
      K3_12882 <= data_out(407 downto 280);
      RConstant_4_12882 <= data_out(279 downto 272);
      K2_12877 <= data_out(271 downto 144);
      RConstant_3_12877 <= data_out(143 downto 136);
      K1_12872 <= data_out(135 downto 8);
      RConstant_2_12872 <= data_out(7 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 1360,
        owidth => 136,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 4,
        nreqs => 10,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => key_expand_single_call_reqs(0),
          ackR => key_expand_single_call_acks(0),
          dataR => key_expand_single_call_data(135 downto 0),
          tagR => key_expand_single_call_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 136,
          owidth => 1360,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 4,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 10) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => key_expand_single_return_acks(0), -- cross-over
          ackL => key_expand_single_return_reqs(0), -- cross-over
          dataL => key_expand_single_return_data(135 downto 0),
          tagL => key_expand_single_return_tag(3 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    call_stmt_12949_call_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= call_stmt_12949_call_req_0;
      call_stmt_12949_call_ack_0<= sample_ack(0);
      update_req(0) <= call_stmt_12949_call_req_1;
      call_stmt_12949_call_ack_1<= update_ack(0);
      call_stmt_12949_call: dec_round_Operator  port map ( -- 
        sample_req => sample_req(0), 
        sample_ack => sample_ack(0), 
        update_req => update_req(0), 
        update_ack => update_ack(0), 
        round_in => round_S10_12941,
        key_in => K9_12940_delayed_1_12944,
        l_round => R_LAST_12947_wire_constant,
        round_out => round_S9_12949,
        clk => clk, reset => reset  
        -- 
      );-- 
    end block;
    call_stmt_12957_call_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= call_stmt_12957_call_req_0;
      call_stmt_12957_call_ack_0<= sample_ack(0);
      update_req(0) <= call_stmt_12957_call_req_1;
      call_stmt_12957_call_ack_1<= update_ack(0);
      call_stmt_12957_call: dec_round_Operator  port map ( -- 
        sample_req => sample_req(0), 
        sample_ack => sample_ack(0), 
        update_req => update_req(0), 
        update_ack => update_ack(0), 
        round_in => round_S9_12949,
        key_in => K8_12945_delayed_2_12952,
        l_round => R_NOT_LAST_12955_wire_constant,
        round_out => round_S8_12957,
        clk => clk, reset => reset  
        -- 
      );-- 
    end block;
    call_stmt_12965_call_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= call_stmt_12965_call_req_0;
      call_stmt_12965_call_ack_0<= sample_ack(0);
      update_req(0) <= call_stmt_12965_call_req_1;
      call_stmt_12965_call_ack_1<= update_ack(0);
      call_stmt_12965_call: dec_round_Operator  port map ( -- 
        sample_req => sample_req(0), 
        sample_ack => sample_ack(0), 
        update_req => update_req(0), 
        update_ack => update_ack(0), 
        round_in => round_S8_12957,
        key_in => K7_12950_delayed_3_12960,
        l_round => R_NOT_LAST_12963_wire_constant,
        round_out => round_S7_12965,
        clk => clk, reset => reset  
        -- 
      );-- 
    end block;
    call_stmt_12973_call_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= call_stmt_12973_call_req_0;
      call_stmt_12973_call_ack_0<= sample_ack(0);
      update_req(0) <= call_stmt_12973_call_req_1;
      call_stmt_12973_call_ack_1<= update_ack(0);
      call_stmt_12973_call: dec_round_Operator  port map ( -- 
        sample_req => sample_req(0), 
        sample_ack => sample_ack(0), 
        update_req => update_req(0), 
        update_ack => update_ack(0), 
        round_in => round_S7_12965,
        key_in => K6_12955_delayed_4_12968,
        l_round => R_NOT_LAST_12971_wire_constant,
        round_out => round_S6_12973,
        clk => clk, reset => reset  
        -- 
      );-- 
    end block;
    call_stmt_12981_call_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= call_stmt_12981_call_req_0;
      call_stmt_12981_call_ack_0<= sample_ack(0);
      update_req(0) <= call_stmt_12981_call_req_1;
      call_stmt_12981_call_ack_1<= update_ack(0);
      call_stmt_12981_call: dec_round_Operator  port map ( -- 
        sample_req => sample_req(0), 
        sample_ack => sample_ack(0), 
        update_req => update_req(0), 
        update_ack => update_ack(0), 
        round_in => round_S6_12973,
        key_in => K5_12960_delayed_5_12976,
        l_round => R_NOT_LAST_12979_wire_constant,
        round_out => round_S5_12981,
        clk => clk, reset => reset  
        -- 
      );-- 
    end block;
    call_stmt_12989_call_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= call_stmt_12989_call_req_0;
      call_stmt_12989_call_ack_0<= sample_ack(0);
      update_req(0) <= call_stmt_12989_call_req_1;
      call_stmt_12989_call_ack_1<= update_ack(0);
      call_stmt_12989_call: dec_round_Operator  port map ( -- 
        sample_req => sample_req(0), 
        sample_ack => sample_ack(0), 
        update_req => update_req(0), 
        update_ack => update_ack(0), 
        round_in => round_S5_12981,
        key_in => K4_12965_delayed_6_12984,
        l_round => R_NOT_LAST_12987_wire_constant,
        round_out => round_S4_12989,
        clk => clk, reset => reset  
        -- 
      );-- 
    end block;
    call_stmt_12997_call_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= call_stmt_12997_call_req_0;
      call_stmt_12997_call_ack_0<= sample_ack(0);
      update_req(0) <= call_stmt_12997_call_req_1;
      call_stmt_12997_call_ack_1<= update_ack(0);
      call_stmt_12997_call: dec_round_Operator  port map ( -- 
        sample_req => sample_req(0), 
        sample_ack => sample_ack(0), 
        update_req => update_req(0), 
        update_ack => update_ack(0), 
        round_in => round_S4_12989,
        key_in => K3_12970_delayed_7_12992,
        l_round => R_NOT_LAST_12995_wire_constant,
        round_out => round_S3_12997,
        clk => clk, reset => reset  
        -- 
      );-- 
    end block;
    call_stmt_13005_call_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= call_stmt_13005_call_req_0;
      call_stmt_13005_call_ack_0<= sample_ack(0);
      update_req(0) <= call_stmt_13005_call_req_1;
      call_stmt_13005_call_ack_1<= update_ack(0);
      call_stmt_13005_call: dec_round_Operator  port map ( -- 
        sample_req => sample_req(0), 
        sample_ack => sample_ack(0), 
        update_req => update_req(0), 
        update_ack => update_ack(0), 
        round_in => round_S3_12997,
        key_in => K2_12975_delayed_8_13000,
        l_round => R_NOT_LAST_13003_wire_constant,
        round_out => round_S2_13005,
        clk => clk, reset => reset  
        -- 
      );-- 
    end block;
    call_stmt_13013_call_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= call_stmt_13013_call_req_0;
      call_stmt_13013_call_ack_0<= sample_ack(0);
      update_req(0) <= call_stmt_13013_call_req_1;
      call_stmt_13013_call_ack_1<= update_ack(0);
      call_stmt_13013_call: dec_round_Operator  port map ( -- 
        sample_req => sample_req(0), 
        sample_ack => sample_ack(0), 
        update_req => update_req(0), 
        update_ack => update_ack(0), 
        round_in => round_S2_13005,
        key_in => K1_12980_delayed_9_13008,
        l_round => R_NOT_LAST_13011_wire_constant,
        round_out => round_S1_13013,
        clk => clk, reset => reset  
        -- 
      );-- 
    end block;
    call_stmt_13021_call_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= call_stmt_13021_call_req_0;
      call_stmt_13021_call_ack_0<= sample_ack(0);
      update_req(0) <= call_stmt_13021_call_req_1;
      call_stmt_13021_call_ack_1<= update_ack(0);
      call_stmt_13021_call: dec_round_Operator  port map ( -- 
        sample_req => sample_req(0), 
        sample_ack => sample_ack(0), 
        update_req => update_req(0), 
        update_ack => update_ack(0), 
        round_in => round_S1_13013,
        key_in => K0_12985_delayed_10_13016,
        l_round => R_NOT_LAST_13019_wire_constant,
        round_out => round_S0_13021,
        clk => clk, reset => reset  
        -- 
      );-- 
    end block;
    -- 
  end Block; -- data_path
  -- 
end d_block_daemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library work;
use work.ahir_system_global_package.all;
entity dec_round_Operator is -- 
  port ( -- 
    sample_req: in boolean;
    sample_ack: out boolean;
    update_req: in boolean;
    update_ack: out boolean;
    round_in : in  std_logic_vector(127 downto 0);
    key_in : in  std_logic_vector(127 downto 0);
    l_round : in  std_logic_vector(0 downto 0);
    round_out : out  std_logic_vector(127 downto 0);
    clk, reset: in std_logic
    -- 
  );
  -- 
end entity dec_round_Operator;
architecture dec_round_Operator_arch of dec_round_Operator is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal update_ack_symbol: Boolean;
  signal default_zero_sig: std_logic;
  -- input port buffer signals
  signal round_in_buffer :  std_logic_vector(127 downto 0);
  signal round_in_update_enable: Boolean;
  signal round_in_update_enable_unmarked: Boolean;
  signal key_in_buffer :  std_logic_vector(127 downto 0);
  signal key_in_update_enable: Boolean;
  signal key_in_update_enable_unmarked: Boolean;
  signal l_round_buffer :  std_logic_vector(0 downto 0);
  signal l_round_update_enable: Boolean;
  signal l_round_update_enable_unmarked: Boolean;
  -- output port buffer signals
  signal round_out_buffer :  std_logic_vector(127 downto 0);
  signal round_out_update_enable: Boolean;
  signal dec_round_CP_3275_start: Boolean;
  signal dec_round_CP_3275_symbol: Boolean;
  signal cp_all_inputs_sampled: Boolean;
  -- volatile/operator module components. 
  component Inv_Sbox_1_Volatile is -- 
    port ( -- 
      s_in : in  std_logic_vector(7 downto 0);
      s_out : out  std_logic_vector(7 downto 0)-- 
    );
    -- 
  end component; 
  component Inv_Sbox_2_Volatile is -- 
    port ( -- 
      s_in : in  std_logic_vector(7 downto 0);
      s_out : out  std_logic_vector(7 downto 0)-- 
    );
    -- 
  end component; 
  component Inv_Sbox_3_Volatile is -- 
    port ( -- 
      s_in : in  std_logic_vector(7 downto 0);
      s_out : out  std_logic_vector(7 downto 0)-- 
    );
    -- 
  end component; 
  component Inv_Sbox_4_Volatile is -- 
    port ( -- 
      s_in : in  std_logic_vector(7 downto 0);
      s_out : out  std_logic_vector(7 downto 0)-- 
    );
    -- 
  end component; 
  component MUL2_Volatile is -- 
    port ( -- 
      mul_in : in  std_logic_vector(7 downto 0);
      mul_out : out  std_logic_vector(7 downto 0)-- 
    );
    -- 
  end component; 
  -- links between control-path and data-path
  signal XOR_u128_u128_12816_inst_req_0 : boolean;
  signal XOR_u128_u128_12816_inst_ack_0 : boolean;
  signal XOR_u128_u128_12816_inst_req_1 : boolean;
  signal XOR_u128_u128_12816_inst_ack_1 : boolean;
  -- 
begin --  
  sample_ack <= dec_round_CP_3275_symbol;
  -- input handling ------------------------------------------------
  round_in_buffer <= round_in;
  key_in_buffer <= key_in;
  l_round_buffer <= l_round;
  dec_round_CP_3275_start <= sample_req;
  -- output handling  -------------------------------------------------------
  round_out <= round_out_buffer;
  round_out_update_enable <= update_req;
  update_ack_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 22) := "update_ack_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= dec_round_CP_3275_symbol & update_req;
    gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => update_ack_symbol, clk => clk, reset => reset); --
  end block;
  -- update ack. 
  update_ack <= update_ack_symbol;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  dec_round_CP_3275: Block -- control-path 
    signal dec_round_CP_3275_elements: BooleanArray(2 downto 0);
    -- 
  begin -- 
    dec_round_CP_3275_elements(0) <= dec_round_CP_3275_start;
    dec_round_CP_3275_symbol <= dec_round_CP_3275_elements(2);
    -- CP-element group 0:  join  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (2852) 
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12162_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12198_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12198_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISa_12189_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12194_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12162_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12162_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12174_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12174_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12162_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12162_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_round_in_12173_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISa_12189_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISa_12189_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12190_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12190_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12198_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12198_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12190_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12194_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12194_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12190_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12186_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12198_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12198_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12186_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISb_12193_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12162_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_round_in_12173_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_round_in_12173_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12162_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_round_in_12173_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12174_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12186_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12186_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12186_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12198_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12198_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12186_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISb_12193_update_start_
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISa_12185_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12174_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_round_in_12161_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_round_in_12161_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12174_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12174_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12186_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12186_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISa_12185_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISb_12197_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISb_12197_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISa_12185_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISb_12193_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISb_12193_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12194_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISa_12185_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12186_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISb_12197_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISb_12197_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12186_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12194_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_round_in_12161_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12170_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12170_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12170_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_round_in_12161_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12170_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12170_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12186_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12186_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12182_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12182_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12198_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12198_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12182_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12194_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12162_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12170_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12170_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12170_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_round_in_12169_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_round_in_12169_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12182_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12182_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12182_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12198_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12198_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12182_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12194_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12190_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12190_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12182_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12194_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12194_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISa_12181_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12190_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_round_in_12169_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_round_in_12169_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12170_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12170_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12170_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12170_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISa_12181_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISa_12181_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISa_12181_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12182_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12194_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12194_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12182_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12190_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12166_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12166_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12166_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12166_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12166_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12182_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12182_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12178_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12178_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12194_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12318_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12178_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12190_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12190_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12178_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12210_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12210_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12178_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12190_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12178_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12178_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12178_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12166_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISa_12177_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISa_12177_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISa_12177_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISa_12177_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12178_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12178_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12190_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12178_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12178_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12202_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12202_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12174_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISa_12189_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12166_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12166_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_round_in_12165_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12174_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12174_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12174_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_round_in_12165_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_round_in_12165_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12174_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_round_in_12165_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12162_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12162_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12166_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12166_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12166_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12166_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12162_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12162_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12174_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12318_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12318_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12202_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12202_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISb_12201_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISb_12201_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISb_12201_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISb_12201_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12202_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12202_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12202_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12202_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12202_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12202_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12202_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12202_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12206_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12206_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12206_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12206_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISb_12205_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISb_12205_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISb_12205_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISb_12205_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12206_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12206_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12206_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12206_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12206_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12206_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12206_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12206_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12210_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12210_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12210_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12210_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISc_12209_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISc_12209_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISc_12209_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISc_12209_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12210_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12210_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12210_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12210_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12263_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12263_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12210_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12210_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12214_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12214_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12214_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12214_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISc_12213_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISc_12213_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISc_12213_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISc_12213_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12214_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12214_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12214_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12214_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12214_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12214_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12214_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12214_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12218_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12218_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12218_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12218_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISc_12217_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISc_12217_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISc_12217_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISc_12217_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12218_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12218_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12218_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12218_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12218_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12218_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12218_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12218_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12486_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12222_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12222_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12222_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12222_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISc_12221_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISc_12221_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISc_12221_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISc_12221_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12486_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS01x2_12485_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12222_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12222_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12222_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12222_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12222_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12222_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12222_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12222_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12492_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12603_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS01x2_12485_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12226_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12226_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12226_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12226_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISd_12225_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISd_12225_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISd_12225_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISd_12225_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_B10_12490_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12226_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12226_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12226_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12226_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12226_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12226_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12226_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12226_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12486_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12486_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS00x2_12484_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS00x2_12484_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12230_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12230_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12230_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12230_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISd_12229_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISd_12229_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISd_12229_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISd_12229_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12496_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12230_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12230_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12487_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12230_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12230_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12230_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12230_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12487_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12230_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12230_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12492_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12492_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12234_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12234_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12234_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12234_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISd_12233_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISd_12233_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISd_12233_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISd_12233_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12234_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12234_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12234_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12234_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12234_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12234_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12234_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12234_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12492_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12496_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12238_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12238_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12238_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12238_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISd_12237_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISd_12237_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISd_12237_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISd_12237_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12238_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12238_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12238_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12238_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12238_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12238_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS00x2_12484_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12238_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/slice_12238_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12242_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12242_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12242_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12242_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS01_12491_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12487_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS00_12240_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS00_12240_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS00_12240_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS00_12240_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12492_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS01x2_12485_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12245_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12245_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12245_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12245_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12487_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS01_12243_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS01_12243_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS01_12243_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS01_12243_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12248_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12248_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12248_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12248_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS00x2_12484_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12486_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS02_12246_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS02_12246_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS02_12246_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS02_12246_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12492_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12487_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12251_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12251_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12251_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12251_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS03_12249_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS03_12249_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS03_12249_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS03_12249_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12496_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12486_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12254_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12254_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12254_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12254_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12486_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12487_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS04_12252_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS04_12252_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS04_12252_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS04_12252_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12486_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12257_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12257_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12257_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12257_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_B10_12490_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS05_12255_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS05_12255_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS05_12255_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS05_12255_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12496_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12260_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12260_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12260_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12260_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS06_12258_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS06_12258_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS06_12258_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS06_12258_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12492_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12492_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12492_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12487_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12263_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS12x2_12340_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS14x2_12341_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS14x2_12341_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS14x2_12341_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS14x2_12341_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12495_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12495_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12263_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12486_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS07_12261_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS07_12261_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS07_12261_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS07_12261_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12266_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12266_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12266_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12266_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS08_12264_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS08_12264_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS08_12264_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS08_12264_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS01_12491_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12269_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12269_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12269_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12269_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12487_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS09_12267_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS09_12267_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS09_12267_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS09_12267_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12492_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12272_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12272_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12272_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12272_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS10_12270_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS10_12270_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS10_12270_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS10_12270_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_B10_12490_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12275_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12275_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12275_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12275_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS01_12491_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS11_12273_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS11_12273_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS11_12273_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS11_12273_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12278_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12278_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12278_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12278_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS12_12276_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS12_12276_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS12_12276_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS12_12276_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12281_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12281_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12281_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12281_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_B10_12490_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12492_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS13_12279_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS13_12279_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS13_12279_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS13_12279_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS01_12491_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12492_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12284_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12284_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12284_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12284_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS14_12282_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS14_12282_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS14_12282_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS14_12282_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS01x2_12485_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12287_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12287_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12287_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12287_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS15_12285_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS15_12285_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS15_12285_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS15_12285_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12295_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12295_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12295_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12295_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12291_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12291_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12291_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12291_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS00_12289_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS00_12289_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS00_12289_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS00_12289_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS01_12290_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS01_12290_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS01_12290_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS01_12290_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12291_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12291_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12291_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12291_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12291_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12291_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12291_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12291_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12294_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12294_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12294_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12294_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS02_12292_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS02_12292_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS02_12292_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS02_12292_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS03_12293_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS03_12293_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS03_12293_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS03_12293_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12294_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12294_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12294_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12294_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12294_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12294_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12294_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12294_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12295_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12295_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12295_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12295_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12295_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12295_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12295_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12295_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12304_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12304_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12304_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12304_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12300_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12300_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12300_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12300_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS04_12298_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS04_12298_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS04_12298_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS04_12298_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS05_12299_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS05_12299_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS05_12299_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS05_12299_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12300_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12300_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12300_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12300_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12300_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12300_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12300_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12300_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12303_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12303_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12303_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12303_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS06_12301_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS06_12301_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS06_12301_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS06_12301_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS07_12302_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS07_12302_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS07_12302_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS07_12302_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12303_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12303_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12303_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12303_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12303_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12303_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12303_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12303_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12304_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12304_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12304_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12304_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12304_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12304_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12304_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12304_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12313_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12313_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12313_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12313_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12309_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12309_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12309_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12309_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS08_12307_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS08_12307_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS08_12307_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS08_12307_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS09_12308_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS09_12308_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS09_12308_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS09_12308_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12309_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12309_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12309_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12309_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12309_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12309_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12309_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12309_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12312_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12312_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12312_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12312_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS10_12310_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS10_12310_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS10_12310_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS10_12310_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS11_12311_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS11_12311_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS11_12311_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS11_12311_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12312_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12312_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12312_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12312_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12312_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12312_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12312_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12312_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12313_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12313_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12313_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12313_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12313_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12313_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12313_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12313_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12322_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12322_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12322_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12322_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12318_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12318_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12318_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12318_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS12_12316_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS12_12316_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS12_12316_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS12_12316_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS13_12317_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS13_12317_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS13_12317_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS13_12317_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12318_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12318_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12318_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12318_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12318_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12321_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12321_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12321_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12321_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS14_12319_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS14_12319_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS14_12319_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS14_12319_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS15_12320_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS15_12320_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS15_12320_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS15_12320_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12321_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12321_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12321_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12321_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12321_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12321_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12321_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12321_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12322_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12322_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12322_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12322_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12322_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12322_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12322_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12322_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12327_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12327_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12327_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12327_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS00x2_12325_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS00x2_12325_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS00x2_12325_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS00x2_12325_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS02x2_12326_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS02x2_12326_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS02x2_12326_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS02x2_12326_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12327_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12327_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12327_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12327_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12327_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12327_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12327_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12327_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12332_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12332_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12332_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12332_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS04x2_12330_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS04x2_12330_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS04x2_12330_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS04x2_12330_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS06x2_12331_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS06x2_12331_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS06x2_12331_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS06x2_12331_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12332_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12332_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12332_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12332_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12332_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12332_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12332_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12332_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12337_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12337_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12337_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12337_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS08x2_12335_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS08x2_12335_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS08x2_12335_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS08x2_12335_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS10x2_12336_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS10x2_12336_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS10x2_12336_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS10x2_12336_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12337_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12337_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12337_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12337_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12337_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12337_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12337_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12337_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12342_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12342_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12342_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12342_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS12x2_12340_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS12x2_12340_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS12x2_12340_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS00x2_12512_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS00x2_12512_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS00x2_12512_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12603_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12600_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12603_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12600_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12603_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12603_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12342_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12342_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12342_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12342_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12342_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12342_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12342_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12342_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12347_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12347_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12347_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12347_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS01x2_12345_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS01x2_12345_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS01x2_12345_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS01x2_12345_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS03x2_12346_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS03x2_12346_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS03x2_12346_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS03x2_12346_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12347_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12347_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12347_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12347_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12347_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12347_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12347_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12347_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12352_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12352_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12352_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12352_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS05x2_12350_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS05x2_12350_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS05x2_12350_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS05x2_12350_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS07x2_12351_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS07x2_12351_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS07x2_12351_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS07x2_12351_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12352_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12352_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12352_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12352_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12352_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12352_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12352_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12352_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12357_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12357_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12357_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12357_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS09x2_12355_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS09x2_12355_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS09x2_12355_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS09x2_12355_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS11x2_12356_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS11x2_12356_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS11x2_12356_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS11x2_12356_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12357_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12357_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12357_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12357_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12357_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12357_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12357_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12357_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12362_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12362_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12362_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12362_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS13x2_12360_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS13x2_12360_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS13x2_12360_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS13x2_12360_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS15x2_12361_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS15x2_12361_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS15x2_12361_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS15x2_12361_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12362_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12362_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12362_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12362_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12362_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12362_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12362_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12362_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12366_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12366_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12366_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12366_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Y00_12364_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Y00_12364_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Y00_12364_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Y00_12364_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12369_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12369_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12369_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12369_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Y01_12367_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Y01_12367_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Y01_12367_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Y01_12367_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12372_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12372_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12372_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12372_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Y02_12370_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Y02_12370_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Y02_12370_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Y02_12370_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12375_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12375_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12375_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12375_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Y03_12373_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Y03_12373_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Y03_12373_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Y03_12373_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12378_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12378_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12378_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12378_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Y10_12376_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Y10_12376_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Y10_12376_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Y10_12376_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12381_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12381_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12381_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12381_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Y11_12379_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Y11_12379_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Y11_12379_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Y11_12379_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12384_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12384_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12384_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12384_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Y12_12382_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Y12_12382_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Y12_12382_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Y12_12382_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12387_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12387_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12387_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12387_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Y13_12385_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Y13_12385_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Y13_12385_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Y13_12385_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12391_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12391_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12391_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12391_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Y00x2_12389_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Y00x2_12389_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Y00x2_12389_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Y00x2_12389_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Y10x2_12390_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Y10x2_12390_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Y10x2_12390_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Y10x2_12390_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12391_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12391_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12391_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12391_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12391_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12391_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12391_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12391_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12600_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12396_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12396_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12396_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12396_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Y01x2_12394_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Y01x2_12394_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Y01x2_12394_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Y01x2_12394_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12604_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12600_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Y11x2_12395_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Y11x2_12395_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Y11x2_12395_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Y11x2_12395_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS14x2_12602_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12396_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12396_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12396_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12396_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12396_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12396_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12396_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12396_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS14_12608_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12603_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12401_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12401_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12401_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12401_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Y02x2_12399_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Y02x2_12399_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Y02x2_12399_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Y02x2_12399_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12613_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12609_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Y12x2_12400_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Y12x2_12400_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Y12x2_12400_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Y12x2_12400_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12609_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12401_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12401_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12401_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12401_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12401_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12401_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12401_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12401_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12406_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12406_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12406_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12406_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Y03x2_12404_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Y03x2_12404_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Y03x2_12404_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Y03x2_12404_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12603_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Y13x2_12405_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Y13x2_12405_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Y13x2_12405_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Y13x2_12405_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12613_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12406_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12406_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12406_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12406_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12406_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12406_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12603_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12406_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12406_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12609_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12609_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS14_12608_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS14_12608_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12410_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12410_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12410_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12410_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12613_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Z0_12408_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Z0_12408_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Z0_12408_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Z0_12408_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12603_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12413_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12413_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12413_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12413_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS14x2_12602_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12609_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Z1_12411_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Z1_12411_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Z1_12411_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Z1_12411_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_B03_12607_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12604_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12416_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12416_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12416_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12416_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Z2_12414_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Z2_12414_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Z2_12414_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Z2_12414_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12419_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12419_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12419_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12419_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12604_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12600_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12609_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Z3_12417_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Z3_12417_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Z3_12417_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Z3_12417_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12609_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12423_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12423_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12423_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12423_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Z0x2_12421_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Z0x2_12421_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Z0x2_12421_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Z0x2_12421_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12600_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12613_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Wc0_12422_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Wc0_12422_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Wc0_12422_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Wc0_12422_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12603_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS13x2_12601_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12604_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12423_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12423_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12423_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12423_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12423_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12423_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12423_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12423_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12609_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u8_u16_12774_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12609_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_B03_12607_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12428_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12428_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12428_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12428_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Z1x2_12426_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Z1x2_12426_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Z1x2_12426_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Z1x2_12426_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_B03_12607_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Wc1_12427_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Wc1_12427_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Wc1_12427_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Wc1_12427_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12428_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12428_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12428_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12428_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12428_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12428_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12428_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12428_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12609_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12433_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12433_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12433_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12433_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Z2x2_12431_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Z2x2_12431_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Z2x2_12431_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Z2x2_12431_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12603_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS13x2_12601_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12604_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Wc2_12432_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Wc2_12432_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Wc2_12432_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Wc2_12432_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_B03_12607_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12609_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12609_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS13x2_12601_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12433_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12433_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12433_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12433_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12433_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12433_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12433_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12433_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS14_12608_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS14x2_12602_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12438_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12438_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12438_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12438_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Z3x2_12436_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Z3x2_12436_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Z3x2_12436_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Z3x2_12436_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12603_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS13x2_12601_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12604_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Wc3_12437_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Wc3_12437_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Wc3_12437_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Wc3_12437_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12438_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12438_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12604_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12438_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12438_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12438_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12438_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12604_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12438_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12438_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS14x2_12602_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12443_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12443_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12443_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12443_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_A0_12441_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_A0_12441_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_A0_12441_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_A0_12441_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Y00x2_12442_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Y00x2_12442_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Y00x2_12442_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Y00x2_12442_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12443_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12443_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12443_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12443_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12443_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12443_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12443_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12443_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12448_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12448_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12448_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12448_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_A1_12446_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_A1_12446_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_A1_12446_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_A1_12446_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Y01x2_12447_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Y01x2_12447_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Y01x2_12447_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Y01x2_12447_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12448_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12448_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12448_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12448_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12448_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12448_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12448_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12448_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12453_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12453_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12453_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12453_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_A2_12451_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_A2_12451_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_A2_12451_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_A2_12451_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Y02x2_12452_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Y02x2_12452_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Y02x2_12452_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Y02x2_12452_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12453_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12453_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12453_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12453_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12453_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12453_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12453_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12453_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12458_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12458_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12458_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12458_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_A3_12456_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_A3_12456_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_A3_12456_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_A3_12456_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Y03x2_12457_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Y03x2_12457_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Y03x2_12457_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Y03x2_12457_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12458_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12458_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12458_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12458_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12458_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12458_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12458_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12458_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12463_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12463_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12463_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12463_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_A0_12461_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_A0_12461_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_A0_12461_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_A0_12461_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Y10x2_12462_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Y10x2_12462_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Y10x2_12462_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Y10x2_12462_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12463_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12463_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12463_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12463_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12463_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12463_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12463_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12463_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12468_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12468_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12468_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12468_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_A1_12466_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_A1_12466_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_A1_12466_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_A1_12466_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Y11x2_12467_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Y11x2_12467_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Y11x2_12467_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Y11x2_12467_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12468_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12468_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12468_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12468_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12468_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12468_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12468_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12468_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12473_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12473_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12473_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12473_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_A2_12471_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_A2_12471_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_A2_12471_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_A2_12471_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Y12x2_12472_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Y12x2_12472_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Y12x2_12472_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Y12x2_12472_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12473_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12473_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12473_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12473_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12473_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12473_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12473_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12473_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12478_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12478_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12478_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12478_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_A3_12476_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_A3_12476_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_A3_12476_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_A3_12476_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Y13x2_12477_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Y13x2_12477_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Y13x2_12477_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Y13x2_12477_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12478_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12478_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12478_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12478_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12478_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12478_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12478_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12478_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12487_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12487_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12487_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12487_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12483_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12483_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12483_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12483_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_B00_12481_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_B00_12481_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_B00_12481_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_B00_12481_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS00_12482_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS00_12482_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS00_12482_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS00_12482_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12483_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12483_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12483_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12483_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12483_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12483_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12483_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12483_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12486_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12486_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12486_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12495_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12495_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS01x2_12493_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS01x2_12493_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS01x2_12493_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS01x2_12493_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS02x2_12494_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS02x2_12494_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS02x2_12494_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS02x2_12494_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12495_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12495_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12495_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12495_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12495_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12495_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12495_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12495_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12496_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12496_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12496_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12496_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12496_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12496_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12496_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12496_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12505_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12505_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12505_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12505_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12501_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12501_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12501_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12501_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_B00_12499_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_B00_12499_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_B00_12499_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_B00_12499_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS02_12500_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS02_12500_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS02_12500_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS02_12500_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12501_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12501_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12501_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12501_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12501_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12501_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12501_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12501_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12504_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12504_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12504_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12504_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS02x2_12502_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS02x2_12502_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS02x2_12502_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS02x2_12502_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS03x2_12503_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS03x2_12503_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS03x2_12503_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS03x2_12503_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12504_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12504_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12504_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12504_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12504_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12504_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12504_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12504_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12505_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12505_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12505_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12505_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12505_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12505_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12505_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12505_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12514_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12514_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12514_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12514_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12510_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12510_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12510_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12510_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_B10_12508_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_B10_12508_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_B10_12508_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_B10_12508_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS03_12509_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS03_12509_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS03_12509_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS03_12509_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12510_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12510_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12510_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12510_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12510_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12510_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12510_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12510_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12513_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12513_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12513_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12513_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS03x2_12511_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS03x2_12511_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS03x2_12511_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS03x2_12511_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS00x2_12512_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12513_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12513_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12513_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12513_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12513_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12513_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12513_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12513_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12514_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12514_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12514_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12514_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12514_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12514_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12514_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12514_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12523_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12523_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12523_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12523_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12519_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12519_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12519_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12519_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_B01_12517_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_B01_12517_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_B01_12517_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_B01_12517_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS04_12518_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS04_12518_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS04_12518_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS04_12518_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12519_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12519_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12519_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12519_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12519_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12519_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12519_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12519_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12522_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12522_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12522_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12522_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS04x2_12520_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS04x2_12520_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS04x2_12520_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS04x2_12520_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS05x2_12521_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS05x2_12521_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS05x2_12521_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS05x2_12521_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12522_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12522_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12522_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12522_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12522_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12522_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12522_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12522_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12523_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12523_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12523_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12523_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12523_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12523_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12523_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12523_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12532_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12532_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12532_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12532_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12528_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12528_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12528_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12528_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_B11_12526_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_B11_12526_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_B11_12526_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_B11_12526_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS05_12527_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS05_12527_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS05_12527_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS05_12527_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12528_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12528_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12528_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12528_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12528_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12528_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12528_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12528_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12531_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12531_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12531_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12531_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS05x2_12529_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS05x2_12529_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS05x2_12529_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS05x2_12529_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS06x2_12530_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS06x2_12530_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS06x2_12530_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS06x2_12530_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12531_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12531_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12531_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12531_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12531_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12531_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12531_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12531_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12532_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12532_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12532_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12532_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12532_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12532_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12532_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12532_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12541_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12541_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12541_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12541_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12537_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12537_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12537_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12537_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_B01_12535_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_B01_12535_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_B01_12535_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_B01_12535_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u8_u16_12771_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u16_u32_12775_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS06_12536_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS06_12536_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS06_12536_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS06_12536_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u16_u32_12784_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12537_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12537_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Sout03_12773_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12537_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12537_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12537_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12537_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u8_u16_12774_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12537_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12537_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u8_u16_12780_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u8_u16_12771_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u8_u16_12774_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u8_u16_12774_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12540_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12540_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12540_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12540_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS06x2_12538_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS06x2_12538_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS06x2_12538_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS06x2_12538_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS07x2_12539_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS07x2_12539_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS07x2_12539_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS07x2_12539_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u8_u16_12774_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u8_u16_12774_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12540_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12540_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12540_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12540_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12540_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12540_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12540_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12540_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u8_u16_12774_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12541_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12541_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u8_u16_12774_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12541_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12541_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12541_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12541_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Sout01_12770_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12541_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12541_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u8_u16_12771_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12550_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12550_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12550_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12550_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12546_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12546_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12546_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12546_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_B11_12544_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_B11_12544_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_B11_12544_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_B11_12544_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS07_12545_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS07_12545_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS07_12545_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS07_12545_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u8_u16_12771_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u16_u32_12784_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Sout00_12769_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12546_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12546_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12546_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12546_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12546_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12546_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12546_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12546_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u8_u16_12774_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12549_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12549_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12549_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12549_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS07x2_12547_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS07x2_12547_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS07x2_12547_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS07x2_12547_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Sout02_12772_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS04x2_12548_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS04x2_12548_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS04x2_12548_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS04x2_12548_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u16_u32_12784_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12549_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12549_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u8_u16_12771_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12549_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12549_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12549_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12549_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u8_u16_12771_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12549_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12549_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u8_u16_12771_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12550_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12550_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12550_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12550_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12550_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12550_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u8_u16_12774_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12550_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12550_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u16_u32_12784_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u16_u32_12775_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12559_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12559_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12559_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12559_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12555_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12555_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12555_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12555_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_B02_12553_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_B02_12553_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_B02_12553_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_B02_12553_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS08_12554_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS08_12554_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS08_12554_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS08_12554_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12555_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12555_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u8_u16_12774_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12555_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12555_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12555_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12555_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12555_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12555_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Sout01_12770_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u16_u32_12775_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u8_u16_12771_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u8_u16_12780_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u16_u32_12775_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Sout02_12772_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12558_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12558_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12558_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12558_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS08x2_12556_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS08x2_12556_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS08x2_12556_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS08x2_12556_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS09x2_12557_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS09x2_12557_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS09x2_12557_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS09x2_12557_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Sout02_12772_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Sout02_12772_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12558_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12558_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u8_u16_12774_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12558_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12558_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12558_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12558_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u16_u32_12775_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12558_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12558_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u8_u16_12780_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u16_u32_12775_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Sout04_12778_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Sout03_12773_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12559_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12559_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Sout01_12770_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12559_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12559_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12559_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12559_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u16_u32_12775_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12559_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12559_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u16_u32_12775_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12568_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12568_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12568_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12568_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12564_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12564_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12564_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12564_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_B12_12562_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_B12_12562_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_B12_12562_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_B12_12562_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Sout01_12770_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Sout04_12778_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS09_12563_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS09_12563_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS09_12563_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS09_12563_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Sout03_12773_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Sout03_12773_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12564_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12564_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12564_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12564_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12564_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12564_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12564_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12564_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u8_u16_12780_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12567_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12567_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12567_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12567_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS09x2_12565_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS09x2_12565_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS09x2_12565_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS09x2_12565_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS10x2_12566_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS10x2_12566_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS10x2_12566_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS10x2_12566_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12567_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12567_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12567_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12567_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12567_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12567_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12567_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12567_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12568_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12568_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12568_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12568_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12568_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12568_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12568_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12568_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12577_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12577_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12577_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12577_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12573_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12573_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12573_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12573_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_B02_12571_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_B02_12571_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_B02_12571_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_B02_12571_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS10_12572_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS10_12572_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS10_12572_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS10_12572_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12573_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12573_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12573_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12573_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12573_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12573_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12573_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12573_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12576_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12576_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12576_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12576_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS10x2_12574_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS10x2_12574_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS10x2_12574_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS10x2_12574_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS11x2_12575_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS11x2_12575_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS11x2_12575_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS11x2_12575_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12576_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12576_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12576_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12576_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12576_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12576_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12576_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12576_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12577_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12577_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12577_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12577_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12577_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12577_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12577_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12577_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12586_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12586_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12586_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12586_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12582_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12582_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12582_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12582_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_B12_12580_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_B12_12580_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_B12_12580_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_B12_12580_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS11_12581_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS11_12581_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS11_12581_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS11_12581_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12582_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12582_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12582_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12582_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12582_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12582_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12582_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12582_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12585_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12585_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12585_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12585_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS11x2_12583_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS11x2_12583_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS11x2_12583_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS11x2_12583_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS08x2_12584_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS08x2_12584_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS08x2_12584_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS08x2_12584_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12585_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12585_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12585_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12585_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12585_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12585_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12585_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12585_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12586_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12586_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12586_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12586_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12586_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12586_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12586_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12586_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12595_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12595_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12595_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12595_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12591_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12591_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12591_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12591_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_B03_12589_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_B03_12589_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_B03_12589_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_B03_12589_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS12_12590_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS12_12590_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS12_12590_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS12_12590_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12591_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12591_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12591_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12591_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12591_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12591_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12591_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12591_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12594_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12594_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12594_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12594_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS12x2_12592_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS12x2_12592_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS12x2_12592_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS12x2_12592_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS13x2_12593_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS13x2_12593_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS13x2_12593_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS13x2_12593_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12594_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12594_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12594_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12594_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12594_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12594_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12594_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12594_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12595_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12595_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12595_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12595_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12595_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12595_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12595_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12595_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12604_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12604_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12604_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12604_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12600_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12600_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12600_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12600_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_B13_12598_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_B13_12598_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_B13_12598_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_B13_12598_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS13_12599_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS13_12599_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS13_12599_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS13_12599_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12600_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12600_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12612_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12612_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12612_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12612_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS14x2_12610_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS14x2_12610_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS14x2_12610_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS14x2_12610_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS15x2_12611_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS15x2_12611_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS15x2_12611_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS15x2_12611_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12612_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12612_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12612_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12612_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12612_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12612_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12612_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12612_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12613_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12613_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12613_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12613_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12613_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12613_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12613_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12613_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12622_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12622_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12622_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12622_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12618_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12618_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12618_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12618_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_B13_12616_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_B13_12616_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_B13_12616_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_B13_12616_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS15_12617_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS15_12617_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS15_12617_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS15_12617_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12618_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12618_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12618_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12618_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12618_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12618_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12618_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12618_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12621_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12621_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12621_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12621_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS15x2_12619_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS15x2_12619_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS15x2_12619_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS15x2_12619_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS12x2_12620_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS12x2_12620_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS12x2_12620_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS12x2_12620_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12621_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12621_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12621_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12621_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12621_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12621_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12621_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12621_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12622_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12622_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12622_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12622_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12622_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12622_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12622_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u8_u8_12622_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12628_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12628_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12628_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12628_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_l_round_12625_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_l_round_12625_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_l_round_12625_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_l_round_12625_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS00_12626_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS00_12626_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS00_12626_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS00_12626_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IMX00_12627_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IMX00_12627_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IMX00_12627_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IMX00_12627_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12628_start/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12628_start/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12628_start/req
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12628_start/ack
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12628_complete/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12628_complete/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12628_complete/req
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12628_complete/ack
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12634_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12634_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12634_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12634_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_l_round_12631_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_l_round_12631_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_l_round_12631_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_l_round_12631_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS01_12632_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS01_12632_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS01_12632_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS01_12632_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IMX01_12633_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IMX01_12633_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IMX01_12633_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IMX01_12633_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12634_start/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12634_start/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12634_start/req
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12634_start/ack
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12634_complete/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12634_complete/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12634_complete/req
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12634_complete/ack
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12640_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12640_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12640_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12640_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_l_round_12637_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_l_round_12637_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_l_round_12637_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_l_round_12637_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS02_12638_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS02_12638_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS02_12638_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS02_12638_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IMX02_12639_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IMX02_12639_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IMX02_12639_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IMX02_12639_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12640_start/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12640_start/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12640_start/req
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12640_start/ack
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12640_complete/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12640_complete/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12640_complete/req
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12640_complete/ack
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12646_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12646_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12646_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12646_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_l_round_12643_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_l_round_12643_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_l_round_12643_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_l_round_12643_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS03_12644_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS03_12644_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS03_12644_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS03_12644_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IMX03_12645_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IMX03_12645_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IMX03_12645_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IMX03_12645_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12646_start/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12646_start/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12646_start/req
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12646_start/ack
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12646_complete/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12646_complete/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12646_complete/req
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12646_complete/ack
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12652_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12652_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12652_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12652_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_l_round_12649_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_l_round_12649_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_l_round_12649_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_l_round_12649_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS04_12650_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS04_12650_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS04_12650_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS04_12650_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IMX04_12651_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IMX04_12651_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IMX04_12651_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IMX04_12651_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12652_start/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12652_start/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12652_start/req
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12652_start/ack
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12652_complete/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12652_complete/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12652_complete/req
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12652_complete/ack
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12658_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12658_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12658_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12658_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_l_round_12655_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_l_round_12655_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_l_round_12655_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_l_round_12655_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS05_12656_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS05_12656_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS05_12656_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS05_12656_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IMX05_12657_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IMX05_12657_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IMX05_12657_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IMX05_12657_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12658_start/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12658_start/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12658_start/req
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12658_start/ack
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12658_complete/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12658_complete/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12658_complete/req
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12658_complete/ack
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12664_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12664_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12664_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12664_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_l_round_12661_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_l_round_12661_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_l_round_12661_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_l_round_12661_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS06_12662_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS06_12662_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS06_12662_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS06_12662_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IMX06_12663_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IMX06_12663_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IMX06_12663_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IMX06_12663_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12664_start/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12664_start/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12664_start/req
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12664_start/ack
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12664_complete/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12664_complete/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12664_complete/req
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12664_complete/ack
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12670_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12670_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12670_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12670_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_l_round_12667_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_l_round_12667_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_l_round_12667_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_l_round_12667_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS07_12668_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS07_12668_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS07_12668_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS07_12668_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IMX07_12669_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IMX07_12669_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IMX07_12669_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IMX07_12669_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12670_start/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12670_start/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12670_start/req
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12670_start/ack
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12670_complete/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12670_complete/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12670_complete/req
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12670_complete/ack
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12676_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12676_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12676_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12676_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_l_round_12673_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_l_round_12673_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_l_round_12673_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_l_round_12673_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS08_12674_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS08_12674_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS08_12674_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS08_12674_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IMX08_12675_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IMX08_12675_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IMX08_12675_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IMX08_12675_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12676_start/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12676_start/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12676_start/req
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12676_start/ack
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12676_complete/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12676_complete/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12676_complete/req
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12676_complete/ack
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12682_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12682_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12682_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12682_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_l_round_12679_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_l_round_12679_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_l_round_12679_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_l_round_12679_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS09_12680_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS09_12680_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS09_12680_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS09_12680_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IMX09_12681_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IMX09_12681_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IMX09_12681_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IMX09_12681_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12682_start/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12682_start/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12682_start/req
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12682_start/ack
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12682_complete/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12682_complete/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12682_complete/req
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12682_complete/ack
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12688_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12688_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12688_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12688_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_l_round_12685_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_l_round_12685_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_l_round_12685_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_l_round_12685_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS10_12686_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS10_12686_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS10_12686_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS10_12686_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IMX10_12687_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IMX10_12687_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IMX10_12687_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IMX10_12687_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12688_start/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12688_start/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12688_start/req
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12688_start/ack
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12688_complete/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12688_complete/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12688_complete/req
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12688_complete/ack
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12694_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12694_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12694_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12694_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_l_round_12691_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_l_round_12691_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_l_round_12691_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_l_round_12691_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS11_12692_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS11_12692_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS11_12692_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS11_12692_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IMX11_12693_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IMX11_12693_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IMX11_12693_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IMX11_12693_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12694_start/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12694_start/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12694_start/req
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12694_start/ack
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12694_complete/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12694_complete/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12694_complete/req
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12694_complete/ack
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12700_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12700_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12700_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12700_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_l_round_12697_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_l_round_12697_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_l_round_12697_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_l_round_12697_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS12_12698_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS12_12698_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS12_12698_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS12_12698_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IMX12_12699_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IMX12_12699_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IMX12_12699_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IMX12_12699_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12700_start/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12700_start/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12700_start/req
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12700_start/ack
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12700_complete/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12700_complete/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12700_complete/req
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12700_complete/ack
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12706_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12706_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12706_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12706_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_l_round_12703_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_l_round_12703_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_l_round_12703_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_l_round_12703_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS13_12704_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS13_12704_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS13_12704_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS13_12704_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IMX13_12705_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IMX13_12705_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IMX13_12705_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IMX13_12705_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12706_start/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12706_start/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12706_start/req
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12706_start/ack
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12706_complete/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12706_complete/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12706_complete/req
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12706_complete/ack
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12712_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12712_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12712_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12712_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_l_round_12709_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_l_round_12709_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_l_round_12709_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_l_round_12709_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS14_12710_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS14_12710_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS14_12710_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS14_12710_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IMX14_12711_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IMX14_12711_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IMX14_12711_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IMX14_12711_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12712_start/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12712_start/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12712_start/req
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12712_start/ack
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12712_complete/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12712_complete/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12712_complete/req
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12712_complete/ack
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12718_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12718_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12718_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12718_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_l_round_12715_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_l_round_12715_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_l_round_12715_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_l_round_12715_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS15_12716_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS15_12716_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS15_12716_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IS15_12716_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IMX15_12717_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IMX15_12717_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IMX15_12717_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_IMX15_12717_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12718_start/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12718_start/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12718_start/req
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12718_start/ack
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12718_complete/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12718_complete/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12718_complete/req
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/MUX_12718_complete/ack
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12722_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12722_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12722_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12722_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISbox_in00_12720_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISbox_in00_12720_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISbox_in00_12720_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISbox_in00_12720_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12725_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12725_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12725_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12725_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISbox_in01_12723_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISbox_in01_12723_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISbox_in01_12723_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISbox_in01_12723_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12728_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12728_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12728_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12728_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISbox_in02_12726_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISbox_in02_12726_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISbox_in02_12726_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISbox_in02_12726_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12731_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12731_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12731_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12731_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISbox_in03_12729_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISbox_in03_12729_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISbox_in03_12729_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISbox_in03_12729_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12734_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12734_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12734_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12734_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISbox_in04_12732_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISbox_in04_12732_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISbox_in04_12732_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISbox_in04_12732_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12737_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12737_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12737_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12737_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISbox_in05_12735_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISbox_in05_12735_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISbox_in05_12735_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISbox_in05_12735_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12740_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12740_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12740_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12740_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISbox_in06_12738_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISbox_in06_12738_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISbox_in06_12738_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISbox_in06_12738_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12743_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12743_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12743_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12743_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISbox_in07_12741_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISbox_in07_12741_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISbox_in07_12741_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISbox_in07_12741_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12746_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12746_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12746_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12746_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISbox_in08_12744_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISbox_in08_12744_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISbox_in08_12744_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISbox_in08_12744_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12749_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12749_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12749_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12749_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISbox_in09_12747_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISbox_in09_12747_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISbox_in09_12747_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISbox_in09_12747_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12752_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12752_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12752_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12752_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISbox_in10_12750_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISbox_in10_12750_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISbox_in10_12750_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISbox_in10_12750_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12755_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12755_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12755_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12755_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISbox_in11_12753_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISbox_in11_12753_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISbox_in11_12753_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISbox_in11_12753_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12758_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12758_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12758_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12758_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISbox_in12_12756_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISbox_in12_12756_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISbox_in12_12756_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISbox_in12_12756_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12761_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12761_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12761_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12761_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISbox_in13_12759_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISbox_in13_12759_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISbox_in13_12759_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISbox_in13_12759_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12764_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12764_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12764_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12764_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISbox_in14_12762_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISbox_in14_12762_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISbox_in14_12762_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISbox_in14_12762_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12767_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12767_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12767_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/call_stmt_12767_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISbox_in15_12765_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISbox_in15_12765_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISbox_in15_12765_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISbox_in15_12765_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u16_u32_12775_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u16_u32_12775_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u16_u32_12775_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u16_u32_12775_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u8_u16_12771_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u8_u16_12771_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u8_u16_12771_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u8_u16_12771_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Sout00_12769_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Sout00_12769_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Sout00_12769_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Sout04_12778_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Sout04_12778_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Sout05_12779_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Sout05_12779_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Sout05_12779_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Sout05_12779_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u8_u16_12780_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u8_u16_12780_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u8_u16_12780_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u8_u16_12780_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u8_u16_12780_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u8_u16_12780_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u8_u16_12780_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u8_u16_12780_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u8_u16_12783_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u8_u16_12783_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u8_u16_12783_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u8_u16_12783_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Sout06_12781_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Sout06_12781_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Sout06_12781_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Sout06_12781_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Sout07_12782_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Sout07_12782_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Sout07_12782_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Sout07_12782_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u8_u16_12783_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u8_u16_12783_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u8_u16_12783_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u8_u16_12783_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u8_u16_12783_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u8_u16_12783_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u8_u16_12783_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u8_u16_12783_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u16_u32_12784_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u16_u32_12784_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u16_u32_12784_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u16_u32_12784_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u16_u32_12784_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u16_u32_12784_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u16_u32_12784_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u16_u32_12784_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u16_u32_12793_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u16_u32_12793_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u16_u32_12793_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u16_u32_12793_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u8_u16_12789_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u8_u16_12789_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u8_u16_12789_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u8_u16_12789_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Sout08_12787_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Sout08_12787_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Sout08_12787_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Sout08_12787_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Sout09_12788_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Sout09_12788_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Sout09_12788_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Sout09_12788_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u8_u16_12789_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u8_u16_12789_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u8_u16_12789_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u8_u16_12789_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u8_u16_12789_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u8_u16_12789_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u8_u16_12789_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u8_u16_12789_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u8_u16_12792_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u8_u16_12792_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u8_u16_12792_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u8_u16_12792_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Sout10_12790_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Sout10_12790_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Sout10_12790_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Sout10_12790_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Sout11_12791_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Sout11_12791_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Sout11_12791_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Sout11_12791_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u8_u16_12792_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u8_u16_12792_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u8_u16_12792_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u8_u16_12792_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u8_u16_12792_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u8_u16_12792_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u8_u16_12792_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u8_u16_12792_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u16_u32_12793_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u16_u32_12793_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u16_u32_12793_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u16_u32_12793_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u16_u32_12793_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u16_u32_12793_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u16_u32_12793_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u16_u32_12793_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u16_u32_12802_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u16_u32_12802_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u16_u32_12802_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u16_u32_12802_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u8_u16_12798_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u8_u16_12798_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u8_u16_12798_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u8_u16_12798_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Sout12_12796_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Sout12_12796_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Sout12_12796_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Sout12_12796_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Sout13_12797_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Sout13_12797_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Sout13_12797_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Sout13_12797_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u8_u16_12798_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u8_u16_12798_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u8_u16_12798_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u8_u16_12798_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u8_u16_12798_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u8_u16_12798_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u8_u16_12798_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u8_u16_12798_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u8_u16_12801_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u8_u16_12801_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u8_u16_12801_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u8_u16_12801_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Sout14_12799_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Sout14_12799_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Sout14_12799_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Sout14_12799_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Sout15_12800_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Sout15_12800_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Sout15_12800_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_Sout15_12800_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u8_u16_12801_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u8_u16_12801_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u8_u16_12801_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u8_u16_12801_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u8_u16_12801_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u8_u16_12801_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u8_u16_12801_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u8_u16_12801_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u16_u32_12802_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u16_u32_12802_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u16_u32_12802_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u16_u32_12802_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u16_u32_12802_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u16_u32_12802_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u16_u32_12802_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u16_u32_12802_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u64_u128_12811_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u64_u128_12811_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u64_u128_12811_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u64_u128_12811_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u32_u64_12807_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u32_u64_12807_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u32_u64_12807_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u32_u64_12807_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISX0_12805_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISX0_12805_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISX0_12805_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISX0_12805_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISX1_12806_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISX1_12806_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISX1_12806_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISX1_12806_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u32_u64_12807_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u32_u64_12807_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u32_u64_12807_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u32_u64_12807_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u32_u64_12807_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u32_u64_12807_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u32_u64_12807_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u32_u64_12807_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u32_u64_12810_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u32_u64_12810_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u32_u64_12810_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u32_u64_12810_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISX2_12808_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISX2_12808_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISX2_12808_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISX2_12808_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISX3_12809_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISX3_12809_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISX3_12809_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_ISX3_12809_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u32_u64_12810_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u32_u64_12810_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u32_u64_12810_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u32_u64_12810_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u32_u64_12810_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u32_u64_12810_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u32_u64_12810_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u32_u64_12810_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u64_u128_12811_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u64_u128_12811_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u64_u128_12811_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u64_u128_12811_Sample/ra
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u64_u128_12811_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u64_u128_12811_Update/$exit
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u64_u128_12811_Update/cr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/CONCAT_u64_u128_12811_Update/ca
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u128_u128_12816_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u128_u128_12816_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_OUT_12814_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_OUT_12814_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_OUT_12814_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_OUT_12814_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_key_in_12815_sample_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_key_in_12815_sample_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_key_in_12815_update_start_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/R_key_in_12815_update_completed_
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u128_u128_12816_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u128_u128_12816_Sample/rr
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u128_u128_12816_Update/$entry
      -- CP-element group 0: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u128_u128_12816_Update/cr
      -- 
    cr_6407_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6407_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dec_round_CP_3275_elements(0), ack => XOR_u128_u128_12816_inst_req_1); -- 
    rr_6402_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6402_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dec_round_CP_3275_elements(0), ack => XOR_u128_u128_12816_inst_req_0); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u128_u128_12816_sample_completed_
      -- CP-element group 1: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u128_u128_12816_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u128_u128_12816_Sample/ra
      -- 
    ra_6403_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => XOR_u128_u128_12816_inst_ack_0, ack => dec_round_CP_3275_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2:  members (5) 
      -- CP-element group 2: 	 assign_stmt_12163_to_assign_stmt_12817/$exit
      -- CP-element group 2: 	 $exit
      -- CP-element group 2: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u128_u128_12816_update_completed_
      -- CP-element group 2: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u128_u128_12816_Update/$exit
      -- CP-element group 2: 	 assign_stmt_12163_to_assign_stmt_12817/XOR_u128_u128_12816_Update/ca
      -- 
    ca_6408_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => XOR_u128_u128_12816_inst_ack_1, ack => dec_round_CP_3275_elements(2)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal A0_12424 : std_logic_vector(7 downto 0);
    signal A1_12429 : std_logic_vector(7 downto 0);
    signal A2_12434 : std_logic_vector(7 downto 0);
    signal A3_12439 : std_logic_vector(7 downto 0);
    signal B00_12444 : std_logic_vector(7 downto 0);
    signal B01_12449 : std_logic_vector(7 downto 0);
    signal B02_12454 : std_logic_vector(7 downto 0);
    signal B03_12459 : std_logic_vector(7 downto 0);
    signal B10_12464 : std_logic_vector(7 downto 0);
    signal B11_12469 : std_logic_vector(7 downto 0);
    signal B12_12474 : std_logic_vector(7 downto 0);
    signal B13_12479 : std_logic_vector(7 downto 0);
    signal CONCAT_u32_u64_12807_wire : std_logic_vector(63 downto 0);
    signal CONCAT_u32_u64_12810_wire : std_logic_vector(63 downto 0);
    signal CONCAT_u8_u16_12771_wire : std_logic_vector(15 downto 0);
    signal CONCAT_u8_u16_12774_wire : std_logic_vector(15 downto 0);
    signal CONCAT_u8_u16_12780_wire : std_logic_vector(15 downto 0);
    signal CONCAT_u8_u16_12783_wire : std_logic_vector(15 downto 0);
    signal CONCAT_u8_u16_12789_wire : std_logic_vector(15 downto 0);
    signal CONCAT_u8_u16_12792_wire : std_logic_vector(15 downto 0);
    signal CONCAT_u8_u16_12798_wire : std_logic_vector(15 downto 0);
    signal CONCAT_u8_u16_12801_wire : std_logic_vector(15 downto 0);
    signal IMX00_12488 : std_logic_vector(7 downto 0);
    signal IMX01_12497 : std_logic_vector(7 downto 0);
    signal IMX02_12506 : std_logic_vector(7 downto 0);
    signal IMX03_12515 : std_logic_vector(7 downto 0);
    signal IMX04_12524 : std_logic_vector(7 downto 0);
    signal IMX05_12533 : std_logic_vector(7 downto 0);
    signal IMX06_12542 : std_logic_vector(7 downto 0);
    signal IMX07_12551 : std_logic_vector(7 downto 0);
    signal IMX08_12560 : std_logic_vector(7 downto 0);
    signal IMX09_12569 : std_logic_vector(7 downto 0);
    signal IMX10_12578 : std_logic_vector(7 downto 0);
    signal IMX11_12587 : std_logic_vector(7 downto 0);
    signal IMX12_12596 : std_logic_vector(7 downto 0);
    signal IMX13_12605 : std_logic_vector(7 downto 0);
    signal IMX14_12614 : std_logic_vector(7 downto 0);
    signal IMX15_12623 : std_logic_vector(7 downto 0);
    signal IS00_12179 : std_logic_vector(7 downto 0);
    signal IS00x2_12242 : std_logic_vector(7 downto 0);
    signal IS01_12183 : std_logic_vector(7 downto 0);
    signal IS01x2_12245 : std_logic_vector(7 downto 0);
    signal IS02_12187 : std_logic_vector(7 downto 0);
    signal IS02x2_12248 : std_logic_vector(7 downto 0);
    signal IS03_12191 : std_logic_vector(7 downto 0);
    signal IS03x2_12251 : std_logic_vector(7 downto 0);
    signal IS04_12195 : std_logic_vector(7 downto 0);
    signal IS04x2_12254 : std_logic_vector(7 downto 0);
    signal IS05_12199 : std_logic_vector(7 downto 0);
    signal IS05x2_12257 : std_logic_vector(7 downto 0);
    signal IS06_12203 : std_logic_vector(7 downto 0);
    signal IS06x2_12260 : std_logic_vector(7 downto 0);
    signal IS07_12207 : std_logic_vector(7 downto 0);
    signal IS07x2_12263 : std_logic_vector(7 downto 0);
    signal IS08_12211 : std_logic_vector(7 downto 0);
    signal IS08x2_12266 : std_logic_vector(7 downto 0);
    signal IS09_12215 : std_logic_vector(7 downto 0);
    signal IS09x2_12269 : std_logic_vector(7 downto 0);
    signal IS10_12219 : std_logic_vector(7 downto 0);
    signal IS10x2_12272 : std_logic_vector(7 downto 0);
    signal IS11_12223 : std_logic_vector(7 downto 0);
    signal IS11x2_12275 : std_logic_vector(7 downto 0);
    signal IS12_12227 : std_logic_vector(7 downto 0);
    signal IS12x2_12278 : std_logic_vector(7 downto 0);
    signal IS13_12231 : std_logic_vector(7 downto 0);
    signal IS13x2_12281 : std_logic_vector(7 downto 0);
    signal IS14_12235 : std_logic_vector(7 downto 0);
    signal IS14x2_12284 : std_logic_vector(7 downto 0);
    signal IS15_12239 : std_logic_vector(7 downto 0);
    signal IS15x2_12287 : std_logic_vector(7 downto 0);
    signal ISX0_12776 : std_logic_vector(31 downto 0);
    signal ISX1_12785 : std_logic_vector(31 downto 0);
    signal ISX2_12794 : std_logic_vector(31 downto 0);
    signal ISX3_12803 : std_logic_vector(31 downto 0);
    signal ISa_12163 : std_logic_vector(31 downto 0);
    signal ISb_12167 : std_logic_vector(31 downto 0);
    signal ISbox_in00_12629 : std_logic_vector(7 downto 0);
    signal ISbox_in01_12635 : std_logic_vector(7 downto 0);
    signal ISbox_in02_12641 : std_logic_vector(7 downto 0);
    signal ISbox_in03_12647 : std_logic_vector(7 downto 0);
    signal ISbox_in04_12653 : std_logic_vector(7 downto 0);
    signal ISbox_in05_12659 : std_logic_vector(7 downto 0);
    signal ISbox_in06_12665 : std_logic_vector(7 downto 0);
    signal ISbox_in07_12671 : std_logic_vector(7 downto 0);
    signal ISbox_in08_12677 : std_logic_vector(7 downto 0);
    signal ISbox_in09_12683 : std_logic_vector(7 downto 0);
    signal ISbox_in10_12689 : std_logic_vector(7 downto 0);
    signal ISbox_in11_12695 : std_logic_vector(7 downto 0);
    signal ISbox_in12_12701 : std_logic_vector(7 downto 0);
    signal ISbox_in13_12707 : std_logic_vector(7 downto 0);
    signal ISbox_in14_12713 : std_logic_vector(7 downto 0);
    signal ISbox_in15_12719 : std_logic_vector(7 downto 0);
    signal ISc_12171 : std_logic_vector(31 downto 0);
    signal ISd_12175 : std_logic_vector(31 downto 0);
    signal OUT_12812 : std_logic_vector(127 downto 0);
    signal Sout00_12722 : std_logic_vector(7 downto 0);
    signal Sout01_12761 : std_logic_vector(7 downto 0);
    signal Sout02_12752 : std_logic_vector(7 downto 0);
    signal Sout03_12743 : std_logic_vector(7 downto 0);
    signal Sout04_12734 : std_logic_vector(7 downto 0);
    signal Sout05_12725 : std_logic_vector(7 downto 0);
    signal Sout06_12764 : std_logic_vector(7 downto 0);
    signal Sout07_12755 : std_logic_vector(7 downto 0);
    signal Sout08_12746 : std_logic_vector(7 downto 0);
    signal Sout09_12737 : std_logic_vector(7 downto 0);
    signal Sout10_12728 : std_logic_vector(7 downto 0);
    signal Sout11_12767 : std_logic_vector(7 downto 0);
    signal Sout12_12758 : std_logic_vector(7 downto 0);
    signal Sout13_12749 : std_logic_vector(7 downto 0);
    signal Sout14_12740 : std_logic_vector(7 downto 0);
    signal Sout15_12731 : std_logic_vector(7 downto 0);
    signal Wc0_12296 : std_logic_vector(7 downto 0);
    signal Wc1_12305 : std_logic_vector(7 downto 0);
    signal Wc2_12314 : std_logic_vector(7 downto 0);
    signal Wc3_12323 : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_12291_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_12294_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_12300_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_12303_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_12309_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_12312_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_12318_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_12321_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_12483_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_12486_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_12492_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_12495_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_12501_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_12504_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_12510_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_12513_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_12519_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_12522_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_12528_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_12531_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_12537_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_12540_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_12546_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_12549_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_12555_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_12558_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_12564_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_12567_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_12573_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_12576_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_12582_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_12585_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_12591_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_12594_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_12600_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_12603_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_12609_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_12612_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_12618_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_12621_wire : std_logic_vector(7 downto 0);
    signal Y00_12328 : std_logic_vector(7 downto 0);
    signal Y00x2_12366 : std_logic_vector(7 downto 0);
    signal Y01_12333 : std_logic_vector(7 downto 0);
    signal Y01x2_12369 : std_logic_vector(7 downto 0);
    signal Y02_12338 : std_logic_vector(7 downto 0);
    signal Y02x2_12372 : std_logic_vector(7 downto 0);
    signal Y03_12343 : std_logic_vector(7 downto 0);
    signal Y03x2_12375 : std_logic_vector(7 downto 0);
    signal Y10_12348 : std_logic_vector(7 downto 0);
    signal Y10x2_12378 : std_logic_vector(7 downto 0);
    signal Y11_12353 : std_logic_vector(7 downto 0);
    signal Y11x2_12381 : std_logic_vector(7 downto 0);
    signal Y12_12358 : std_logic_vector(7 downto 0);
    signal Y12x2_12384 : std_logic_vector(7 downto 0);
    signal Y13_12363 : std_logic_vector(7 downto 0);
    signal Y13x2_12387 : std_logic_vector(7 downto 0);
    signal Z0_12392 : std_logic_vector(7 downto 0);
    signal Z0x2_12410 : std_logic_vector(7 downto 0);
    signal Z1_12397 : std_logic_vector(7 downto 0);
    signal Z1x2_12413 : std_logic_vector(7 downto 0);
    signal Z2_12402 : std_logic_vector(7 downto 0);
    signal Z2x2_12416 : std_logic_vector(7 downto 0);
    signal Z3_12407 : std_logic_vector(7 downto 0);
    signal Z3x2_12419 : std_logic_vector(7 downto 0);
    signal xxdec_roundxxsel : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    xxdec_roundxxsel <= "01111111";
    -- flow-through select operator MUX_12628_inst
    ISbox_in00_12629 <= IS00_12179 when (l_round_buffer(0) /=  '0') else IMX00_12488;
    -- flow-through select operator MUX_12634_inst
    ISbox_in01_12635 <= IS01_12183 when (l_round_buffer(0) /=  '0') else IMX01_12497;
    -- flow-through select operator MUX_12640_inst
    ISbox_in02_12641 <= IS02_12187 when (l_round_buffer(0) /=  '0') else IMX02_12506;
    -- flow-through select operator MUX_12646_inst
    ISbox_in03_12647 <= IS03_12191 when (l_round_buffer(0) /=  '0') else IMX03_12515;
    -- flow-through select operator MUX_12652_inst
    ISbox_in04_12653 <= IS04_12195 when (l_round_buffer(0) /=  '0') else IMX04_12524;
    -- flow-through select operator MUX_12658_inst
    ISbox_in05_12659 <= IS05_12199 when (l_round_buffer(0) /=  '0') else IMX05_12533;
    -- flow-through select operator MUX_12664_inst
    ISbox_in06_12665 <= IS06_12203 when (l_round_buffer(0) /=  '0') else IMX06_12542;
    -- flow-through select operator MUX_12670_inst
    ISbox_in07_12671 <= IS07_12207 when (l_round_buffer(0) /=  '0') else IMX07_12551;
    -- flow-through select operator MUX_12676_inst
    ISbox_in08_12677 <= IS08_12211 when (l_round_buffer(0) /=  '0') else IMX08_12560;
    -- flow-through select operator MUX_12682_inst
    ISbox_in09_12683 <= IS09_12215 when (l_round_buffer(0) /=  '0') else IMX09_12569;
    -- flow-through select operator MUX_12688_inst
    ISbox_in10_12689 <= IS10_12219 when (l_round_buffer(0) /=  '0') else IMX10_12578;
    -- flow-through select operator MUX_12694_inst
    ISbox_in11_12695 <= IS11_12223 when (l_round_buffer(0) /=  '0') else IMX11_12587;
    -- flow-through select operator MUX_12700_inst
    ISbox_in12_12701 <= IS12_12227 when (l_round_buffer(0) /=  '0') else IMX12_12596;
    -- flow-through select operator MUX_12706_inst
    ISbox_in13_12707 <= IS13_12231 when (l_round_buffer(0) /=  '0') else IMX13_12605;
    -- flow-through select operator MUX_12712_inst
    ISbox_in14_12713 <= IS14_12235 when (l_round_buffer(0) /=  '0') else IMX14_12614;
    -- flow-through select operator MUX_12718_inst
    ISbox_in15_12719 <= IS15_12239 when (l_round_buffer(0) /=  '0') else IMX15_12623;
    -- flow-through slice operator slice_12162_inst
    ISa_12163 <= round_in_buffer(127 downto 96);
    -- flow-through slice operator slice_12166_inst
    ISb_12167 <= round_in_buffer(95 downto 64);
    -- flow-through slice operator slice_12170_inst
    ISc_12171 <= round_in_buffer(63 downto 32);
    -- flow-through slice operator slice_12174_inst
    ISd_12175 <= round_in_buffer(31 downto 0);
    -- flow-through slice operator slice_12178_inst
    IS00_12179 <= ISa_12163(31 downto 24);
    -- flow-through slice operator slice_12182_inst
    IS01_12183 <= ISa_12163(23 downto 16);
    -- flow-through slice operator slice_12186_inst
    IS02_12187 <= ISa_12163(15 downto 8);
    -- flow-through slice operator slice_12190_inst
    IS03_12191 <= ISa_12163(7 downto 0);
    -- flow-through slice operator slice_12194_inst
    IS04_12195 <= ISb_12167(31 downto 24);
    -- flow-through slice operator slice_12198_inst
    IS05_12199 <= ISb_12167(23 downto 16);
    -- flow-through slice operator slice_12202_inst
    IS06_12203 <= ISb_12167(15 downto 8);
    -- flow-through slice operator slice_12206_inst
    IS07_12207 <= ISb_12167(7 downto 0);
    -- flow-through slice operator slice_12210_inst
    IS08_12211 <= ISc_12171(31 downto 24);
    -- flow-through slice operator slice_12214_inst
    IS09_12215 <= ISc_12171(23 downto 16);
    -- flow-through slice operator slice_12218_inst
    IS10_12219 <= ISc_12171(15 downto 8);
    -- flow-through slice operator slice_12222_inst
    IS11_12223 <= ISc_12171(7 downto 0);
    -- flow-through slice operator slice_12226_inst
    IS12_12227 <= ISd_12175(31 downto 24);
    -- flow-through slice operator slice_12230_inst
    IS13_12231 <= ISd_12175(23 downto 16);
    -- flow-through slice operator slice_12234_inst
    IS14_12235 <= ISd_12175(15 downto 8);
    -- flow-through slice operator slice_12238_inst
    IS15_12239 <= ISd_12175(7 downto 0);
    -- binary operator CONCAT_u16_u32_12775_inst
    process(CONCAT_u8_u16_12771_wire, CONCAT_u8_u16_12774_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u8_u16_12771_wire, CONCAT_u8_u16_12774_wire, tmp_var);
      ISX0_12776 <= tmp_var; -- 
    end process;
    -- binary operator CONCAT_u16_u32_12784_inst
    process(CONCAT_u8_u16_12780_wire, CONCAT_u8_u16_12783_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u8_u16_12780_wire, CONCAT_u8_u16_12783_wire, tmp_var);
      ISX1_12785 <= tmp_var; -- 
    end process;
    -- binary operator CONCAT_u16_u32_12793_inst
    process(CONCAT_u8_u16_12789_wire, CONCAT_u8_u16_12792_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u8_u16_12789_wire, CONCAT_u8_u16_12792_wire, tmp_var);
      ISX2_12794 <= tmp_var; -- 
    end process;
    -- binary operator CONCAT_u16_u32_12802_inst
    process(CONCAT_u8_u16_12798_wire, CONCAT_u8_u16_12801_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u8_u16_12798_wire, CONCAT_u8_u16_12801_wire, tmp_var);
      ISX3_12803 <= tmp_var; -- 
    end process;
    -- binary operator CONCAT_u32_u64_12807_inst
    process(ISX0_12776, ISX1_12785) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApConcat_proc(ISX0_12776, ISX1_12785, tmp_var);
      CONCAT_u32_u64_12807_wire <= tmp_var; -- 
    end process;
    -- binary operator CONCAT_u32_u64_12810_inst
    process(ISX2_12794, ISX3_12803) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApConcat_proc(ISX2_12794, ISX3_12803, tmp_var);
      CONCAT_u32_u64_12810_wire <= tmp_var; -- 
    end process;
    -- binary operator CONCAT_u64_u128_12811_inst
    process(CONCAT_u32_u64_12807_wire, CONCAT_u32_u64_12810_wire) -- 
      variable tmp_var : std_logic_vector(127 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u32_u64_12807_wire, CONCAT_u32_u64_12810_wire, tmp_var);
      OUT_12812 <= tmp_var; -- 
    end process;
    -- binary operator CONCAT_u8_u16_12771_inst
    process(Sout00_12722, Sout01_12761) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApConcat_proc(Sout00_12722, Sout01_12761, tmp_var);
      CONCAT_u8_u16_12771_wire <= tmp_var; -- 
    end process;
    -- binary operator CONCAT_u8_u16_12774_inst
    process(Sout02_12752, Sout03_12743) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApConcat_proc(Sout02_12752, Sout03_12743, tmp_var);
      CONCAT_u8_u16_12774_wire <= tmp_var; -- 
    end process;
    -- binary operator CONCAT_u8_u16_12780_inst
    process(Sout04_12734, Sout05_12725) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApConcat_proc(Sout04_12734, Sout05_12725, tmp_var);
      CONCAT_u8_u16_12780_wire <= tmp_var; -- 
    end process;
    -- binary operator CONCAT_u8_u16_12783_inst
    process(Sout06_12764, Sout07_12755) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApConcat_proc(Sout06_12764, Sout07_12755, tmp_var);
      CONCAT_u8_u16_12783_wire <= tmp_var; -- 
    end process;
    -- binary operator CONCAT_u8_u16_12789_inst
    process(Sout08_12746, Sout09_12737) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApConcat_proc(Sout08_12746, Sout09_12737, tmp_var);
      CONCAT_u8_u16_12789_wire <= tmp_var; -- 
    end process;
    -- binary operator CONCAT_u8_u16_12792_inst
    process(Sout10_12728, Sout11_12767) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApConcat_proc(Sout10_12728, Sout11_12767, tmp_var);
      CONCAT_u8_u16_12792_wire <= tmp_var; -- 
    end process;
    -- binary operator CONCAT_u8_u16_12798_inst
    process(Sout12_12758, Sout13_12749) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApConcat_proc(Sout12_12758, Sout13_12749, tmp_var);
      CONCAT_u8_u16_12798_wire <= tmp_var; -- 
    end process;
    -- binary operator CONCAT_u8_u16_12801_inst
    process(Sout14_12740, Sout15_12731) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApConcat_proc(Sout14_12740, Sout15_12731, tmp_var);
      CONCAT_u8_u16_12801_wire <= tmp_var; -- 
    end process;
    -- shared split operator group (15) : XOR_u128_u128_12816_inst 
    ApIntXor_group_15: Block -- 
      signal data_in: std_logic_vector(255 downto 0);
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= OUT_12812 & key_in_buffer;
      round_out_buffer <= data_out(127 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= XOR_u128_u128_12816_inst_req_0;
      XOR_u128_u128_12816_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= XOR_u128_u128_12816_inst_req_1;
      XOR_u128_u128_12816_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(name => "gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntXor",
          name => "ApIntXor_group_15",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 128,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 128, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 128,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 15
    -- binary operator XOR_u8_u8_12291_inst
    process(IS00_12179, IS01_12183) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(IS00_12179, IS01_12183, tmp_var);
      XOR_u8_u8_12291_wire <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_12294_inst
    process(IS02_12187, IS03_12191) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(IS02_12187, IS03_12191, tmp_var);
      XOR_u8_u8_12294_wire <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_12295_inst
    process(XOR_u8_u8_12291_wire, XOR_u8_u8_12294_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(XOR_u8_u8_12291_wire, XOR_u8_u8_12294_wire, tmp_var);
      Wc0_12296 <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_12300_inst
    process(IS04_12195, IS05_12199) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(IS04_12195, IS05_12199, tmp_var);
      XOR_u8_u8_12300_wire <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_12303_inst
    process(IS06_12203, IS07_12207) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(IS06_12203, IS07_12207, tmp_var);
      XOR_u8_u8_12303_wire <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_12304_inst
    process(XOR_u8_u8_12300_wire, XOR_u8_u8_12303_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(XOR_u8_u8_12300_wire, XOR_u8_u8_12303_wire, tmp_var);
      Wc1_12305 <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_12309_inst
    process(IS08_12211, IS09_12215) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(IS08_12211, IS09_12215, tmp_var);
      XOR_u8_u8_12309_wire <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_12312_inst
    process(IS10_12219, IS11_12223) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(IS10_12219, IS11_12223, tmp_var);
      XOR_u8_u8_12312_wire <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_12313_inst
    process(XOR_u8_u8_12309_wire, XOR_u8_u8_12312_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(XOR_u8_u8_12309_wire, XOR_u8_u8_12312_wire, tmp_var);
      Wc2_12314 <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_12318_inst
    process(IS12_12227, IS13_12231) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(IS12_12227, IS13_12231, tmp_var);
      XOR_u8_u8_12318_wire <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_12321_inst
    process(IS14_12235, IS15_12239) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(IS14_12235, IS15_12239, tmp_var);
      XOR_u8_u8_12321_wire <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_12322_inst
    process(XOR_u8_u8_12318_wire, XOR_u8_u8_12321_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(XOR_u8_u8_12318_wire, XOR_u8_u8_12321_wire, tmp_var);
      Wc3_12323 <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_12327_inst
    process(IS00x2_12242, IS02x2_12248) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(IS00x2_12242, IS02x2_12248, tmp_var);
      Y00_12328 <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_12332_inst
    process(IS04x2_12254, IS06x2_12260) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(IS04x2_12254, IS06x2_12260, tmp_var);
      Y01_12333 <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_12337_inst
    process(IS08x2_12266, IS10x2_12272) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(IS08x2_12266, IS10x2_12272, tmp_var);
      Y02_12338 <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_12342_inst
    process(IS12x2_12278, IS14x2_12284) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(IS12x2_12278, IS14x2_12284, tmp_var);
      Y03_12343 <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_12347_inst
    process(IS01x2_12245, IS03x2_12251) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(IS01x2_12245, IS03x2_12251, tmp_var);
      Y10_12348 <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_12352_inst
    process(IS05x2_12257, IS07x2_12263) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(IS05x2_12257, IS07x2_12263, tmp_var);
      Y11_12353 <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_12357_inst
    process(IS09x2_12269, IS11x2_12275) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(IS09x2_12269, IS11x2_12275, tmp_var);
      Y12_12358 <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_12362_inst
    process(IS13x2_12281, IS15x2_12287) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(IS13x2_12281, IS15x2_12287, tmp_var);
      Y13_12363 <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_12391_inst
    process(Y00x2_12366, Y10x2_12378) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(Y00x2_12366, Y10x2_12378, tmp_var);
      Z0_12392 <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_12396_inst
    process(Y01x2_12369, Y11x2_12381) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(Y01x2_12369, Y11x2_12381, tmp_var);
      Z1_12397 <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_12401_inst
    process(Y02x2_12372, Y12x2_12384) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(Y02x2_12372, Y12x2_12384, tmp_var);
      Z2_12402 <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_12406_inst
    process(Y03x2_12375, Y13x2_12387) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(Y03x2_12375, Y13x2_12387, tmp_var);
      Z3_12407 <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_12423_inst
    process(Z0x2_12410, Wc0_12296) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(Z0x2_12410, Wc0_12296, tmp_var);
      A0_12424 <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_12428_inst
    process(Z1x2_12413, Wc1_12305) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(Z1x2_12413, Wc1_12305, tmp_var);
      A1_12429 <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_12433_inst
    process(Z2x2_12416, Wc2_12314) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(Z2x2_12416, Wc2_12314, tmp_var);
      A2_12434 <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_12438_inst
    process(Z3x2_12419, Wc3_12323) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(Z3x2_12419, Wc3_12323, tmp_var);
      A3_12439 <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_12443_inst
    process(A0_12424, Y00x2_12366) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(A0_12424, Y00x2_12366, tmp_var);
      B00_12444 <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_12448_inst
    process(A1_12429, Y01x2_12369) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(A1_12429, Y01x2_12369, tmp_var);
      B01_12449 <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_12453_inst
    process(A2_12434, Y02x2_12372) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(A2_12434, Y02x2_12372, tmp_var);
      B02_12454 <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_12458_inst
    process(A3_12439, Y03x2_12375) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(A3_12439, Y03x2_12375, tmp_var);
      B03_12459 <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_12463_inst
    process(A0_12424, Y10x2_12378) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(A0_12424, Y10x2_12378, tmp_var);
      B10_12464 <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_12468_inst
    process(A1_12429, Y11x2_12381) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(A1_12429, Y11x2_12381, tmp_var);
      B11_12469 <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_12473_inst
    process(A2_12434, Y12x2_12384) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(A2_12434, Y12x2_12384, tmp_var);
      B12_12474 <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_12478_inst
    process(A3_12439, Y13x2_12387) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(A3_12439, Y13x2_12387, tmp_var);
      B13_12479 <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_12483_inst
    process(B00_12444, IS00_12179) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(B00_12444, IS00_12179, tmp_var);
      XOR_u8_u8_12483_wire <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_12486_inst
    process(IS00x2_12242, IS01x2_12245) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(IS00x2_12242, IS01x2_12245, tmp_var);
      XOR_u8_u8_12486_wire <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_12487_inst
    process(XOR_u8_u8_12483_wire, XOR_u8_u8_12486_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(XOR_u8_u8_12483_wire, XOR_u8_u8_12486_wire, tmp_var);
      IMX00_12488 <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_12492_inst
    process(B10_12464, IS01_12183) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(B10_12464, IS01_12183, tmp_var);
      XOR_u8_u8_12492_wire <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_12495_inst
    process(IS01x2_12245, IS02x2_12248) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(IS01x2_12245, IS02x2_12248, tmp_var);
      XOR_u8_u8_12495_wire <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_12496_inst
    process(XOR_u8_u8_12492_wire, XOR_u8_u8_12495_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(XOR_u8_u8_12492_wire, XOR_u8_u8_12495_wire, tmp_var);
      IMX01_12497 <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_12501_inst
    process(B00_12444, IS02_12187) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(B00_12444, IS02_12187, tmp_var);
      XOR_u8_u8_12501_wire <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_12504_inst
    process(IS02x2_12248, IS03x2_12251) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(IS02x2_12248, IS03x2_12251, tmp_var);
      XOR_u8_u8_12504_wire <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_12505_inst
    process(XOR_u8_u8_12501_wire, XOR_u8_u8_12504_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(XOR_u8_u8_12501_wire, XOR_u8_u8_12504_wire, tmp_var);
      IMX02_12506 <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_12510_inst
    process(B10_12464, IS03_12191) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(B10_12464, IS03_12191, tmp_var);
      XOR_u8_u8_12510_wire <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_12513_inst
    process(IS03x2_12251, IS00x2_12242) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(IS03x2_12251, IS00x2_12242, tmp_var);
      XOR_u8_u8_12513_wire <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_12514_inst
    process(XOR_u8_u8_12510_wire, XOR_u8_u8_12513_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(XOR_u8_u8_12510_wire, XOR_u8_u8_12513_wire, tmp_var);
      IMX03_12515 <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_12519_inst
    process(B01_12449, IS04_12195) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(B01_12449, IS04_12195, tmp_var);
      XOR_u8_u8_12519_wire <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_12522_inst
    process(IS04x2_12254, IS05x2_12257) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(IS04x2_12254, IS05x2_12257, tmp_var);
      XOR_u8_u8_12522_wire <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_12523_inst
    process(XOR_u8_u8_12519_wire, XOR_u8_u8_12522_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(XOR_u8_u8_12519_wire, XOR_u8_u8_12522_wire, tmp_var);
      IMX04_12524 <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_12528_inst
    process(B11_12469, IS05_12199) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(B11_12469, IS05_12199, tmp_var);
      XOR_u8_u8_12528_wire <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_12531_inst
    process(IS05x2_12257, IS06x2_12260) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(IS05x2_12257, IS06x2_12260, tmp_var);
      XOR_u8_u8_12531_wire <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_12532_inst
    process(XOR_u8_u8_12528_wire, XOR_u8_u8_12531_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(XOR_u8_u8_12528_wire, XOR_u8_u8_12531_wire, tmp_var);
      IMX05_12533 <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_12537_inst
    process(B01_12449, IS06_12203) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(B01_12449, IS06_12203, tmp_var);
      XOR_u8_u8_12537_wire <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_12540_inst
    process(IS06x2_12260, IS07x2_12263) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(IS06x2_12260, IS07x2_12263, tmp_var);
      XOR_u8_u8_12540_wire <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_12541_inst
    process(XOR_u8_u8_12537_wire, XOR_u8_u8_12540_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(XOR_u8_u8_12537_wire, XOR_u8_u8_12540_wire, tmp_var);
      IMX06_12542 <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_12546_inst
    process(B11_12469, IS07_12207) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(B11_12469, IS07_12207, tmp_var);
      XOR_u8_u8_12546_wire <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_12549_inst
    process(IS07x2_12263, IS04x2_12254) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(IS07x2_12263, IS04x2_12254, tmp_var);
      XOR_u8_u8_12549_wire <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_12550_inst
    process(XOR_u8_u8_12546_wire, XOR_u8_u8_12549_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(XOR_u8_u8_12546_wire, XOR_u8_u8_12549_wire, tmp_var);
      IMX07_12551 <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_12555_inst
    process(B02_12454, IS08_12211) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(B02_12454, IS08_12211, tmp_var);
      XOR_u8_u8_12555_wire <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_12558_inst
    process(IS08x2_12266, IS09x2_12269) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(IS08x2_12266, IS09x2_12269, tmp_var);
      XOR_u8_u8_12558_wire <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_12559_inst
    process(XOR_u8_u8_12555_wire, XOR_u8_u8_12558_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(XOR_u8_u8_12555_wire, XOR_u8_u8_12558_wire, tmp_var);
      IMX08_12560 <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_12564_inst
    process(B12_12474, IS09_12215) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(B12_12474, IS09_12215, tmp_var);
      XOR_u8_u8_12564_wire <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_12567_inst
    process(IS09x2_12269, IS10x2_12272) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(IS09x2_12269, IS10x2_12272, tmp_var);
      XOR_u8_u8_12567_wire <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_12568_inst
    process(XOR_u8_u8_12564_wire, XOR_u8_u8_12567_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(XOR_u8_u8_12564_wire, XOR_u8_u8_12567_wire, tmp_var);
      IMX09_12569 <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_12573_inst
    process(B02_12454, IS10_12219) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(B02_12454, IS10_12219, tmp_var);
      XOR_u8_u8_12573_wire <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_12576_inst
    process(IS10x2_12272, IS11x2_12275) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(IS10x2_12272, IS11x2_12275, tmp_var);
      XOR_u8_u8_12576_wire <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_12577_inst
    process(XOR_u8_u8_12573_wire, XOR_u8_u8_12576_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(XOR_u8_u8_12573_wire, XOR_u8_u8_12576_wire, tmp_var);
      IMX10_12578 <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_12582_inst
    process(B12_12474, IS11_12223) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(B12_12474, IS11_12223, tmp_var);
      XOR_u8_u8_12582_wire <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_12585_inst
    process(IS11x2_12275, IS08x2_12266) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(IS11x2_12275, IS08x2_12266, tmp_var);
      XOR_u8_u8_12585_wire <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_12586_inst
    process(XOR_u8_u8_12582_wire, XOR_u8_u8_12585_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(XOR_u8_u8_12582_wire, XOR_u8_u8_12585_wire, tmp_var);
      IMX11_12587 <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_12591_inst
    process(B03_12459, IS12_12227) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(B03_12459, IS12_12227, tmp_var);
      XOR_u8_u8_12591_wire <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_12594_inst
    process(IS12x2_12278, IS13x2_12281) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(IS12x2_12278, IS13x2_12281, tmp_var);
      XOR_u8_u8_12594_wire <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_12595_inst
    process(XOR_u8_u8_12591_wire, XOR_u8_u8_12594_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(XOR_u8_u8_12591_wire, XOR_u8_u8_12594_wire, tmp_var);
      IMX12_12596 <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_12600_inst
    process(B13_12479, IS13_12231) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(B13_12479, IS13_12231, tmp_var);
      XOR_u8_u8_12600_wire <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_12603_inst
    process(IS13x2_12281, IS14x2_12284) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(IS13x2_12281, IS14x2_12284, tmp_var);
      XOR_u8_u8_12603_wire <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_12604_inst
    process(XOR_u8_u8_12600_wire, XOR_u8_u8_12603_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(XOR_u8_u8_12600_wire, XOR_u8_u8_12603_wire, tmp_var);
      IMX13_12605 <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_12609_inst
    process(B03_12459, IS14_12235) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(B03_12459, IS14_12235, tmp_var);
      XOR_u8_u8_12609_wire <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_12612_inst
    process(IS14x2_12284, IS15x2_12287) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(IS14x2_12284, IS15x2_12287, tmp_var);
      XOR_u8_u8_12612_wire <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_12613_inst
    process(XOR_u8_u8_12609_wire, XOR_u8_u8_12612_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(XOR_u8_u8_12609_wire, XOR_u8_u8_12612_wire, tmp_var);
      IMX14_12614 <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_12618_inst
    process(B13_12479, IS15_12239) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(B13_12479, IS15_12239, tmp_var);
      XOR_u8_u8_12618_wire <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_12621_inst
    process(IS15x2_12287, IS12x2_12278) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(IS15x2_12287, IS12x2_12278, tmp_var);
      XOR_u8_u8_12621_wire <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_12622_inst
    process(XOR_u8_u8_12618_wire, XOR_u8_u8_12621_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(XOR_u8_u8_12618_wire, XOR_u8_u8_12621_wire, tmp_var);
      IMX15_12623 <= tmp_var; -- 
    end process;
    call_inst_17283: MUL2_Volatile port map(mul_in => IS00_12179, mul_out => IS00x2_12242); 
    call_inst_17284: MUL2_Volatile port map(mul_in => IS01_12183, mul_out => IS01x2_12245); 
    call_inst_17285: MUL2_Volatile port map(mul_in => IS02_12187, mul_out => IS02x2_12248); 
    call_inst_17286: MUL2_Volatile port map(mul_in => IS03_12191, mul_out => IS03x2_12251); 
    call_inst_17287: MUL2_Volatile port map(mul_in => IS04_12195, mul_out => IS04x2_12254); 
    call_inst_17288: MUL2_Volatile port map(mul_in => IS05_12199, mul_out => IS05x2_12257); 
    call_inst_17289: MUL2_Volatile port map(mul_in => IS06_12203, mul_out => IS06x2_12260); 
    call_inst_17290: MUL2_Volatile port map(mul_in => IS07_12207, mul_out => IS07x2_12263); 
    call_inst_17291: MUL2_Volatile port map(mul_in => IS08_12211, mul_out => IS08x2_12266); 
    call_inst_17292: MUL2_Volatile port map(mul_in => IS09_12215, mul_out => IS09x2_12269); 
    call_inst_17293: MUL2_Volatile port map(mul_in => IS10_12219, mul_out => IS10x2_12272); 
    call_inst_17294: MUL2_Volatile port map(mul_in => IS11_12223, mul_out => IS11x2_12275); 
    call_inst_17295: MUL2_Volatile port map(mul_in => IS12_12227, mul_out => IS12x2_12278); 
    call_inst_17296: MUL2_Volatile port map(mul_in => IS13_12231, mul_out => IS13x2_12281); 
    call_inst_17297: MUL2_Volatile port map(mul_in => IS14_12235, mul_out => IS14x2_12284); 
    call_inst_17298: MUL2_Volatile port map(mul_in => IS15_12239, mul_out => IS15x2_12287); 
    call_inst_17319: MUL2_Volatile port map(mul_in => Y00_12328, mul_out => Y00x2_12366); 
    call_inst_17320: MUL2_Volatile port map(mul_in => Y01_12333, mul_out => Y01x2_12369); 
    call_inst_17321: MUL2_Volatile port map(mul_in => Y02_12338, mul_out => Y02x2_12372); 
    call_inst_17322: MUL2_Volatile port map(mul_in => Y03_12343, mul_out => Y03x2_12375); 
    call_inst_17323: MUL2_Volatile port map(mul_in => Y10_12348, mul_out => Y10x2_12378); 
    call_inst_17324: MUL2_Volatile port map(mul_in => Y11_12353, mul_out => Y11x2_12381); 
    call_inst_17325: MUL2_Volatile port map(mul_in => Y12_12358, mul_out => Y12x2_12384); 
    call_inst_17326: MUL2_Volatile port map(mul_in => Y13_12363, mul_out => Y13x2_12387); 
    call_inst_17331: MUL2_Volatile port map(mul_in => Z0_12392, mul_out => Z0x2_12410); 
    call_inst_17332: MUL2_Volatile port map(mul_in => Z1_12397, mul_out => Z1x2_12413); 
    call_inst_17333: MUL2_Volatile port map(mul_in => Z2_12402, mul_out => Z2x2_12416); 
    call_inst_17334: MUL2_Volatile port map(mul_in => Z3_12407, mul_out => Z3x2_12419); 
    call_inst_17411: Inv_Sbox_1_Volatile port map(s_in => ISbox_in00_12629, s_out => Sout00_12722); 
    call_inst_17412: Inv_Sbox_2_Volatile port map(s_in => ISbox_in01_12635, s_out => Sout05_12725); 
    call_inst_17413: Inv_Sbox_3_Volatile port map(s_in => ISbox_in02_12641, s_out => Sout10_12728); 
    call_inst_17414: Inv_Sbox_4_Volatile port map(s_in => ISbox_in03_12647, s_out => Sout15_12731); 
    call_inst_17415: Inv_Sbox_1_Volatile port map(s_in => ISbox_in04_12653, s_out => Sout04_12734); 
    call_inst_17416: Inv_Sbox_2_Volatile port map(s_in => ISbox_in05_12659, s_out => Sout09_12737); 
    call_inst_17417: Inv_Sbox_3_Volatile port map(s_in => ISbox_in06_12665, s_out => Sout14_12740); 
    call_inst_17418: Inv_Sbox_4_Volatile port map(s_in => ISbox_in07_12671, s_out => Sout03_12743); 
    call_inst_17419: Inv_Sbox_1_Volatile port map(s_in => ISbox_in08_12677, s_out => Sout08_12746); 
    call_inst_17420: Inv_Sbox_2_Volatile port map(s_in => ISbox_in09_12683, s_out => Sout13_12749); 
    call_inst_17421: Inv_Sbox_3_Volatile port map(s_in => ISbox_in10_12689, s_out => Sout02_12752); 
    call_inst_17422: Inv_Sbox_4_Volatile port map(s_in => ISbox_in11_12695, s_out => Sout07_12755); 
    call_inst_17423: Inv_Sbox_1_Volatile port map(s_in => ISbox_in12_12701, s_out => Sout12_12758); 
    call_inst_17424: Inv_Sbox_2_Volatile port map(s_in => ISbox_in13_12707, s_out => Sout01_12761); 
    call_inst_17425: Inv_Sbox_3_Volatile port map(s_in => ISbox_in14_12713, s_out => Sout06_12764); 
    call_inst_17426: Inv_Sbox_4_Volatile port map(s_in => ISbox_in15_12719, s_out => Sout11_12767); 
    -- 
  end Block; -- data_path
  -- 
end dec_round_Operator_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library work;
use work.ahir_system_global_package.all;
entity e_block_daemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    e_in_buf_pipe_read_req : out  std_logic_vector(0 downto 0);
    e_in_buf_pipe_read_ack : in   std_logic_vector(0 downto 0);
    e_in_buf_pipe_read_data : in   std_logic_vector(127 downto 0);
    e_cmd_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    e_cmd_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    e_cmd_pipe_pipe_read_data : in   std_logic_vector(143 downto 0);
    e_out_buf_pipe_write_req : out  std_logic_vector(0 downto 0);
    e_out_buf_pipe_write_ack : in   std_logic_vector(0 downto 0);
    e_out_buf_pipe_write_data : out  std_logic_vector(127 downto 0);
    e_block_done_pipe_write_req : out  std_logic_vector(0 downto 0);
    e_block_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
    e_block_done_pipe_write_data : out  std_logic_vector(0 downto 0);
    key_expand_single_call_reqs : out  std_logic_vector(0 downto 0);
    key_expand_single_call_acks : in   std_logic_vector(0 downto 0);
    key_expand_single_call_data : out  std_logic_vector(135 downto 0);
    key_expand_single_call_tag  :  out  std_logic_vector(3 downto 0);
    key_expand_single_return_reqs : out  std_logic_vector(0 downto 0);
    key_expand_single_return_acks : in   std_logic_vector(0 downto 0);
    key_expand_single_return_data : in   std_logic_vector(135 downto 0);
    key_expand_single_return_tag :  in   std_logic_vector(3 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity e_block_daemon;
architecture e_block_daemon_arch of e_block_daemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal e_block_daemon_CP_11105_start: Boolean;
  signal e_block_daemon_CP_11105_symbol: Boolean;
  -- volatile/operator module components. 
  component key_expand_single is -- 
    generic (tag_length : integer); 
    port ( -- 
      K_in : in  std_logic_vector(127 downto 0);
      Round_C : in  std_logic_vector(7 downto 0);
      K_out : out  std_logic_vector(127 downto 0);
      nRound_C : out  std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component enc_round_Operator is -- 
    port ( -- 
      sample_req: in boolean;
      sample_ack: out boolean;
      update_req: in boolean;
      update_ack: out boolean;
      round_in : in  std_logic_vector(127 downto 0);
      key_in : in  std_logic_vector(127 downto 0);
      l_round : in  std_logic_vector(0 downto 0);
      round_out : out  std_logic_vector(127 downto 0);
      clk, reset: in std_logic
      -- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal WPIPE_e_block_done_13737_inst_req_1 : boolean;
  signal WPIPE_e_block_done_13737_inst_ack_0 : boolean;
  signal WPIPE_e_block_done_13737_inst_req_0 : boolean;
  signal call_stmt_13811_call_ack_1 : boolean;
  signal WPIPE_e_block_done_13737_inst_ack_1 : boolean;
  signal call_stmt_13811_call_req_1 : boolean;
  signal n_count_var_13933_13833_buf_req_0 : boolean;
  signal phi_stmt_13830_req_0 : boolean;
  signal W_round_S0_13810_delayed_1_13843_inst_ack_1 : boolean;
  signal W_round_S0_13810_delayed_1_13843_inst_req_0 : boolean;
  signal W_round_S0_13810_delayed_1_13843_inst_req_1 : boolean;
  signal RPIPE_e_in_buf_13836_inst_req_1 : boolean;
  signal phi_stmt_13830_ack_0 : boolean;
  signal call_stmt_13816_call_req_0 : boolean;
  signal call_stmt_13816_call_req_1 : boolean;
  signal call_stmt_13816_call_ack_0 : boolean;
  signal call_stmt_13816_call_ack_1 : boolean;
  signal n_count_var_13933_13833_buf_ack_0 : boolean;
  signal RPIPE_e_cmd_pipe_13742_inst_req_0 : boolean;
  signal RPIPE_e_cmd_pipe_13742_inst_ack_0 : boolean;
  signal RPIPE_e_cmd_pipe_13742_inst_req_1 : boolean;
  signal RPIPE_e_cmd_pipe_13742_inst_ack_1 : boolean;
  signal do_while_stmt_13828_branch_req_0 : boolean;
  signal RPIPE_e_in_buf_13836_inst_ack_0 : boolean;
  signal RPIPE_e_in_buf_13836_inst_req_0 : boolean;
  signal W_round_S0_13810_delayed_1_13843_inst_ack_0 : boolean;
  signal call_stmt_13811_call_ack_0 : boolean;
  signal call_stmt_13821_call_ack_1 : boolean;
  signal call_stmt_13821_call_req_1 : boolean;
  signal call_stmt_13811_call_req_0 : boolean;
  signal call_stmt_13821_call_ack_0 : boolean;
  signal call_stmt_13821_call_req_0 : boolean;
  signal if_stmt_13756_branch_req_0 : boolean;
  signal if_stmt_13756_branch_ack_1 : boolean;
  signal if_stmt_13756_branch_ack_0 : boolean;
  signal n_count_var_13933_13833_buf_ack_1 : boolean;
  signal n_count_var_13933_13833_buf_req_1 : boolean;
  signal call_stmt_13776_call_req_0 : boolean;
  signal call_stmt_13776_call_ack_0 : boolean;
  signal call_stmt_13776_call_req_1 : boolean;
  signal call_stmt_13776_call_ack_1 : boolean;
  signal phi_stmt_13830_req_1 : boolean;
  signal call_stmt_13781_call_req_0 : boolean;
  signal call_stmt_13781_call_ack_0 : boolean;
  signal call_stmt_13781_call_req_1 : boolean;
  signal call_stmt_13781_call_ack_1 : boolean;
  signal RPIPE_e_in_buf_13836_inst_ack_1 : boolean;
  signal call_stmt_13786_call_req_0 : boolean;
  signal call_stmt_13786_call_ack_0 : boolean;
  signal call_stmt_13786_call_req_1 : boolean;
  signal call_stmt_13786_call_ack_1 : boolean;
  signal e_new_key_13955_13766_buf_req_1 : boolean;
  signal call_stmt_13791_call_req_0 : boolean;
  signal call_stmt_13791_call_ack_0 : boolean;
  signal call_stmt_13791_call_req_1 : boolean;
  signal call_stmt_13791_call_ack_1 : boolean;
  signal phi_stmt_13763_req_0 : boolean;
  signal call_stmt_13796_call_req_0 : boolean;
  signal call_stmt_13796_call_ack_0 : boolean;
  signal call_stmt_13796_call_req_1 : boolean;
  signal call_stmt_13796_call_ack_1 : boolean;
  signal e_init_key_13755_13765_buf_req_1 : boolean;
  signal call_stmt_13801_call_req_0 : boolean;
  signal call_stmt_13801_call_ack_0 : boolean;
  signal call_stmt_13801_call_req_1 : boolean;
  signal call_stmt_13801_call_ack_1 : boolean;
  signal call_stmt_13806_call_req_0 : boolean;
  signal call_stmt_13806_call_ack_0 : boolean;
  signal call_stmt_13806_call_req_1 : boolean;
  signal call_stmt_13806_call_ack_1 : boolean;
  signal W_K1_13811_delayed_1_13846_inst_req_0 : boolean;
  signal W_K1_13811_delayed_1_13846_inst_ack_0 : boolean;
  signal W_K1_13811_delayed_1_13846_inst_req_1 : boolean;
  signal W_K1_13811_delayed_1_13846_inst_ack_1 : boolean;
  signal call_stmt_13853_call_req_0 : boolean;
  signal call_stmt_13853_call_ack_0 : boolean;
  signal call_stmt_13853_call_req_1 : boolean;
  signal call_stmt_13853_call_ack_1 : boolean;
  signal W_K2_13816_delayed_2_13854_inst_req_0 : boolean;
  signal W_K2_13816_delayed_2_13854_inst_ack_0 : boolean;
  signal W_K2_13816_delayed_2_13854_inst_req_1 : boolean;
  signal W_K2_13816_delayed_2_13854_inst_ack_1 : boolean;
  signal call_stmt_13861_call_req_0 : boolean;
  signal call_stmt_13861_call_ack_0 : boolean;
  signal call_stmt_13861_call_req_1 : boolean;
  signal call_stmt_13861_call_ack_1 : boolean;
  signal W_K3_13821_delayed_3_13862_inst_req_0 : boolean;
  signal W_K3_13821_delayed_3_13862_inst_ack_0 : boolean;
  signal W_K3_13821_delayed_3_13862_inst_req_1 : boolean;
  signal W_K3_13821_delayed_3_13862_inst_ack_1 : boolean;
  signal call_stmt_13869_call_req_0 : boolean;
  signal call_stmt_13869_call_ack_0 : boolean;
  signal call_stmt_13869_call_req_1 : boolean;
  signal call_stmt_13869_call_ack_1 : boolean;
  signal W_K4_13826_delayed_4_13870_inst_req_0 : boolean;
  signal W_K4_13826_delayed_4_13870_inst_ack_0 : boolean;
  signal W_K4_13826_delayed_4_13870_inst_req_1 : boolean;
  signal W_K4_13826_delayed_4_13870_inst_ack_1 : boolean;
  signal call_stmt_13877_call_req_0 : boolean;
  signal call_stmt_13877_call_ack_0 : boolean;
  signal call_stmt_13877_call_req_1 : boolean;
  signal call_stmt_13877_call_ack_1 : boolean;
  signal W_K5_13831_delayed_5_13878_inst_req_0 : boolean;
  signal W_K5_13831_delayed_5_13878_inst_ack_0 : boolean;
  signal W_K5_13831_delayed_5_13878_inst_req_1 : boolean;
  signal W_K5_13831_delayed_5_13878_inst_ack_1 : boolean;
  signal call_stmt_13885_call_req_0 : boolean;
  signal call_stmt_13885_call_ack_0 : boolean;
  signal call_stmt_13885_call_req_1 : boolean;
  signal call_stmt_13885_call_ack_1 : boolean;
  signal W_K6_13836_delayed_6_13886_inst_req_0 : boolean;
  signal W_K6_13836_delayed_6_13886_inst_ack_0 : boolean;
  signal W_K6_13836_delayed_6_13886_inst_req_1 : boolean;
  signal W_K6_13836_delayed_6_13886_inst_ack_1 : boolean;
  signal e_init_key_13755_13765_buf_ack_1 : boolean;
  signal e_init_key_13755_13765_buf_ack_0 : boolean;
  signal call_stmt_13893_call_req_0 : boolean;
  signal call_stmt_13893_call_ack_0 : boolean;
  signal if_stmt_13956_branch_ack_0 : boolean;
  signal call_stmt_13893_call_req_1 : boolean;
  signal call_stmt_13893_call_ack_1 : boolean;
  signal W_K7_13841_delayed_7_13894_inst_req_0 : boolean;
  signal W_K7_13841_delayed_7_13894_inst_ack_0 : boolean;
  signal W_K7_13841_delayed_7_13894_inst_req_1 : boolean;
  signal W_K7_13841_delayed_7_13894_inst_ack_1 : boolean;
  signal e_init_key_13755_13765_buf_req_0 : boolean;
  signal phi_stmt_13767_req_0 : boolean;
  signal e_init_count_13751_13769_buf_ack_1 : boolean;
  signal e_init_count_13751_13769_buf_req_1 : boolean;
  signal e_new_key_13955_13766_buf_ack_0 : boolean;
  signal e_new_key_13955_13766_buf_req_0 : boolean;
  signal if_stmt_13956_branch_ack_1 : boolean;
  signal call_stmt_13901_call_req_0 : boolean;
  signal call_stmt_13901_call_ack_0 : boolean;
  signal call_stmt_13901_call_req_1 : boolean;
  signal call_stmt_13901_call_ack_1 : boolean;
  signal phi_stmt_13767_ack_0 : boolean;
  signal e_new_count_13951_13770_buf_req_0 : boolean;
  signal e_new_count_13951_13770_buf_ack_0 : boolean;
  signal if_stmt_13956_branch_req_0 : boolean;
  signal W_K8_13846_delayed_8_13902_inst_req_0 : boolean;
  signal W_K8_13846_delayed_8_13902_inst_ack_0 : boolean;
  signal W_K8_13846_delayed_8_13902_inst_req_1 : boolean;
  signal W_K8_13846_delayed_8_13902_inst_ack_1 : boolean;
  signal phi_stmt_13763_ack_0 : boolean;
  signal e_init_count_13751_13769_buf_ack_0 : boolean;
  signal call_stmt_13909_call_req_0 : boolean;
  signal call_stmt_13909_call_ack_0 : boolean;
  signal call_stmt_13909_call_req_1 : boolean;
  signal call_stmt_13909_call_ack_1 : boolean;
  signal e_init_count_13751_13769_buf_req_0 : boolean;
  signal W_K9_13851_delayed_9_13910_inst_req_0 : boolean;
  signal W_K9_13851_delayed_9_13910_inst_ack_0 : boolean;
  signal W_K9_13851_delayed_9_13910_inst_req_1 : boolean;
  signal W_K9_13851_delayed_9_13910_inst_ack_1 : boolean;
  signal phi_stmt_13767_req_1 : boolean;
  signal call_stmt_13917_call_req_0 : boolean;
  signal call_stmt_13917_call_ack_0 : boolean;
  signal call_stmt_13917_call_req_1 : boolean;
  signal call_stmt_13917_call_ack_1 : boolean;
  signal e_new_count_13951_13770_buf_req_1 : boolean;
  signal e_new_count_13951_13770_buf_ack_1 : boolean;
  signal W_K10_13856_delayed_10_13918_inst_req_0 : boolean;
  signal W_K10_13856_delayed_10_13918_inst_ack_0 : boolean;
  signal W_K10_13856_delayed_10_13918_inst_req_1 : boolean;
  signal W_K10_13856_delayed_10_13918_inst_ack_1 : boolean;
  signal e_new_key_13955_13766_buf_ack_1 : boolean;
  signal phi_stmt_13763_req_1 : boolean;
  signal call_stmt_13925_call_req_0 : boolean;
  signal call_stmt_13925_call_ack_0 : boolean;
  signal call_stmt_13925_call_req_1 : boolean;
  signal call_stmt_13925_call_ack_1 : boolean;
  signal WPIPE_e_out_buf_13926_inst_req_0 : boolean;
  signal WPIPE_e_out_buf_13926_inst_ack_0 : boolean;
  signal WPIPE_e_out_buf_13926_inst_req_1 : boolean;
  signal WPIPE_e_out_buf_13926_inst_ack_1 : boolean;
  signal ADD_u15_u15_13932_inst_req_0 : boolean;
  signal ADD_u15_u15_13932_inst_ack_0 : boolean;
  signal ADD_u15_u15_13932_inst_req_1 : boolean;
  signal ADD_u15_u15_13932_inst_ack_1 : boolean;
  signal do_while_stmt_13828_branch_ack_0 : boolean;
  signal do_while_stmt_13828_branch_ack_1 : boolean;
  signal WPIPE_e_block_done_13938_inst_req_0 : boolean;
  signal WPIPE_e_block_done_13938_inst_ack_0 : boolean;
  signal WPIPE_e_block_done_13938_inst_req_1 : boolean;
  signal WPIPE_e_block_done_13938_inst_ack_1 : boolean;
  signal RPIPE_e_cmd_pipe_13942_inst_req_0 : boolean;
  signal RPIPE_e_cmd_pipe_13942_inst_ack_0 : boolean;
  signal RPIPE_e_cmd_pipe_13942_inst_req_1 : boolean;
  signal RPIPE_e_cmd_pipe_13942_inst_ack_1 : boolean;
  signal countA_13767_13825_buf_req_0 : boolean;
  signal countA_13767_13825_buf_ack_0 : boolean;
  signal countA_13767_13825_buf_req_1 : boolean;
  signal countA_13767_13825_buf_ack_1 : boolean;
  signal phi_stmt_13823_req_0 : boolean;
  signal e_new_count_13951_13826_buf_req_0 : boolean;
  signal e_new_count_13951_13826_buf_ack_0 : boolean;
  signal e_new_count_13951_13826_buf_req_1 : boolean;
  signal e_new_count_13951_13826_buf_ack_1 : boolean;
  signal phi_stmt_13823_req_1 : boolean;
  signal phi_stmt_13823_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "e_block_daemon_input_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      bypass_flag => true,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  e_block_daemon_CP_11105_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "e_block_daemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= e_block_daemon_CP_11105_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= e_block_daemon_CP_11105_start & tag_ilock_write_ack_symbol;
    gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= e_block_daemon_CP_11105_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  e_block_daemon_CP_11105: Block -- control-path 
    signal e_block_daemon_CP_11105_elements: BooleanArray(249 downto 0);
    -- 
  begin -- 
    e_block_daemon_CP_11105_elements(0) <= e_block_daemon_CP_11105_start;
    -- unreachable exit of control-path
    e_block_daemon_CP_11105_symbol <= false;
    -- CP-element group 0:  transition  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (2) 
      -- CP-element group 0: 	 branch_block_stmt_13736/$entry
      -- CP-element group 0: 	 $entry
      -- 
    -- CP-element group 1:  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	14 
    -- CP-element group 1:  members (2) 
      -- CP-element group 1: 	 branch_block_stmt_13736/assign_stmt_13739__entry__
      -- CP-element group 1: 	 branch_block_stmt_13736/branch_block_stmt_13736__entry__
      -- 
    e_block_daemon_CP_11105_elements(1) <= e_block_daemon_CP_11105_elements(0);
    -- CP-element group 2:  branch  place  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	16 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	210 
    -- CP-element group 2: 	211 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_13736/merge_stmt_13740__entry__
      -- CP-element group 2: 	 branch_block_stmt_13736/assign_stmt_13739__exit__
      -- 
    e_block_daemon_CP_11105_elements(2) <= e_block_daemon_CP_11105_elements(16);
    -- CP-element group 3:  merge  place  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	214 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	17 
    -- CP-element group 3:  members (2) 
      -- CP-element group 3: 	 branch_block_stmt_13736/assign_stmt_13743__entry__
      -- CP-element group 3: 	 branch_block_stmt_13736/merge_stmt_13740__exit__
      -- 
    e_block_daemon_CP_11105_elements(3) <= e_block_daemon_CP_11105_elements(214);
    -- CP-element group 4:  place  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	19 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	20 
    -- CP-element group 4:  members (2) 
      -- CP-element group 4: 	 branch_block_stmt_13736/assign_stmt_13747_to_assign_stmt_13755__entry__
      -- CP-element group 4: 	 branch_block_stmt_13736/assign_stmt_13743__exit__
      -- 
    e_block_daemon_CP_11105_elements(4) <= e_block_daemon_CP_11105_elements(19);
    -- CP-element group 5:  branch  place  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	20 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	21 
    -- CP-element group 5: 	22 
    -- CP-element group 5:  members (2) 
      -- CP-element group 5: 	 branch_block_stmt_13736/if_stmt_13756__entry__
      -- CP-element group 5: 	 branch_block_stmt_13736/assign_stmt_13747_to_assign_stmt_13755__exit__
      -- 
    e_block_daemon_CP_11105_elements(5) <= e_block_daemon_CP_11105_elements(20);
    -- CP-element group 6:  merge  branch  place  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	27 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	215 
    -- CP-element group 6: 	216 
    -- CP-element group 6:  members (2) 
      -- CP-element group 6: 	 branch_block_stmt_13736/merge_stmt_13762__entry__
      -- CP-element group 6: 	 branch_block_stmt_13736/if_stmt_13756__exit__
      -- 
    e_block_daemon_CP_11105_elements(6) <= e_block_daemon_CP_11105_elements(27);
    -- CP-element group 7:  merge  place  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	236 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	29 
    -- CP-element group 7:  members (2) 
      -- CP-element group 7: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821__entry__
      -- CP-element group 7: 	 branch_block_stmt_13736/merge_stmt_13762__exit__
      -- 
    e_block_daemon_CP_11105_elements(7) <= e_block_daemon_CP_11105_elements(236);
    -- CP-element group 8:  branch  place  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	49 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	237 
    -- CP-element group 8: 	238 
    -- CP-element group 8:  members (2) 
      -- CP-element group 8: 	 branch_block_stmt_13736/merge_stmt_13822__entry__
      -- CP-element group 8: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821__exit__
      -- 
    e_block_daemon_CP_11105_elements(8) <= e_block_daemon_CP_11105_elements(49);
    -- CP-element group 9:  merge  place  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	248 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	50 
    -- CP-element group 9:  members (2) 
      -- CP-element group 9: 	 branch_block_stmt_13736/do_while_stmt_13828__entry__
      -- CP-element group 9: 	 branch_block_stmt_13736/merge_stmt_13822__exit__
      -- 
    e_block_daemon_CP_11105_elements(9) <= e_block_daemon_CP_11105_elements(248);
    -- CP-element group 10:  place  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	193 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	194 
    -- CP-element group 10:  members (2) 
      -- CP-element group 10: 	 branch_block_stmt_13736/assign_stmt_13940__entry__
      -- CP-element group 10: 	 branch_block_stmt_13736/do_while_stmt_13828__exit__
      -- 
    e_block_daemon_CP_11105_elements(10) <= e_block_daemon_CP_11105_elements(193);
    -- CP-element group 11:  place  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	196 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	197 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_13736/assign_stmt_13940__exit__
      -- CP-element group 11: 	 branch_block_stmt_13736/assign_stmt_13943__entry__
      -- 
    e_block_daemon_CP_11105_elements(11) <= e_block_daemon_CP_11105_elements(196);
    -- CP-element group 12:  place  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	199 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	200 
    -- CP-element group 12:  members (2) 
      -- CP-element group 12: 	 branch_block_stmt_13736/assign_stmt_13947_to_assign_stmt_13955__entry__
      -- CP-element group 12: 	 branch_block_stmt_13736/assign_stmt_13943__exit__
      -- 
    e_block_daemon_CP_11105_elements(12) <= e_block_daemon_CP_11105_elements(199);
    -- CP-element group 13:  branch  place  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	200 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	201 
    -- CP-element group 13: 	202 
    -- CP-element group 13:  members (2) 
      -- CP-element group 13: 	 branch_block_stmt_13736/if_stmt_13956__entry__
      -- CP-element group 13: 	 branch_block_stmt_13736/assign_stmt_13947_to_assign_stmt_13955__exit__
      -- 
    e_block_daemon_CP_11105_elements(13) <= e_block_daemon_CP_11105_elements(200);
    -- CP-element group 14:  transition  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	1 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (4) 
      -- CP-element group 14: 	 branch_block_stmt_13736/assign_stmt_13739/WPIPE_e_block_done_13737_Sample/req
      -- CP-element group 14: 	 branch_block_stmt_13736/assign_stmt_13739/WPIPE_e_block_done_13737_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_13736/assign_stmt_13739/WPIPE_e_block_done_13737_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_13736/assign_stmt_13739/$entry
      -- 
    req_11149_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_11149_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_block_daemon_CP_11105_elements(14), ack => WPIPE_e_block_done_13737_inst_req_0); -- 
    e_block_daemon_CP_11105_elements(14) <= e_block_daemon_CP_11105_elements(1);
    -- CP-element group 15:  transition  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (6) 
      -- CP-element group 15: 	 branch_block_stmt_13736/assign_stmt_13739/WPIPE_e_block_done_13737_Update/req
      -- CP-element group 15: 	 branch_block_stmt_13736/assign_stmt_13739/WPIPE_e_block_done_13737_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_13736/assign_stmt_13739/WPIPE_e_block_done_13737_Sample/ack
      -- CP-element group 15: 	 branch_block_stmt_13736/assign_stmt_13739/WPIPE_e_block_done_13737_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_13736/assign_stmt_13739/WPIPE_e_block_done_13737_update_start_
      -- CP-element group 15: 	 branch_block_stmt_13736/assign_stmt_13739/WPIPE_e_block_done_13737_sample_completed_
      -- 
    ack_11150_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_e_block_done_13737_inst_ack_0, ack => e_block_daemon_CP_11105_elements(15)); -- 
    req_11154_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_11154_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_block_daemon_CP_11105_elements(15), ack => WPIPE_e_block_done_13737_inst_req_1); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	2 
    -- CP-element group 16:  members (4) 
      -- CP-element group 16: 	 branch_block_stmt_13736/assign_stmt_13739/WPIPE_e_block_done_13737_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_13736/assign_stmt_13739/WPIPE_e_block_done_13737_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_13736/assign_stmt_13739/$exit
      -- CP-element group 16: 	 branch_block_stmt_13736/assign_stmt_13739/WPIPE_e_block_done_13737_Update/ack
      -- 
    ack_11155_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_e_block_done_13737_inst_ack_1, ack => e_block_daemon_CP_11105_elements(16)); -- 
    -- CP-element group 17:  transition  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	3 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (4) 
      -- CP-element group 17: 	 branch_block_stmt_13736/assign_stmt_13743/$entry
      -- CP-element group 17: 	 branch_block_stmt_13736/assign_stmt_13743/RPIPE_e_cmd_pipe_13742_sample_start_
      -- CP-element group 17: 	 branch_block_stmt_13736/assign_stmt_13743/RPIPE_e_cmd_pipe_13742_Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_13736/assign_stmt_13743/RPIPE_e_cmd_pipe_13742_Sample/rr
      -- 
    rr_11166_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11166_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_block_daemon_CP_11105_elements(17), ack => RPIPE_e_cmd_pipe_13742_inst_req_0); -- 
    e_block_daemon_CP_11105_elements(17) <= e_block_daemon_CP_11105_elements(3);
    -- CP-element group 18:  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (6) 
      -- CP-element group 18: 	 branch_block_stmt_13736/assign_stmt_13743/RPIPE_e_cmd_pipe_13742_sample_completed_
      -- CP-element group 18: 	 branch_block_stmt_13736/assign_stmt_13743/RPIPE_e_cmd_pipe_13742_update_start_
      -- CP-element group 18: 	 branch_block_stmt_13736/assign_stmt_13743/RPIPE_e_cmd_pipe_13742_Sample/$exit
      -- CP-element group 18: 	 branch_block_stmt_13736/assign_stmt_13743/RPIPE_e_cmd_pipe_13742_Sample/ra
      -- CP-element group 18: 	 branch_block_stmt_13736/assign_stmt_13743/RPIPE_e_cmd_pipe_13742_Update/$entry
      -- CP-element group 18: 	 branch_block_stmt_13736/assign_stmt_13743/RPIPE_e_cmd_pipe_13742_Update/cr
      -- 
    ra_11167_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_e_cmd_pipe_13742_inst_ack_0, ack => e_block_daemon_CP_11105_elements(18)); -- 
    cr_11171_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11171_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_block_daemon_CP_11105_elements(18), ack => RPIPE_e_cmd_pipe_13742_inst_req_1); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	4 
    -- CP-element group 19:  members (4) 
      -- CP-element group 19: 	 branch_block_stmt_13736/assign_stmt_13743/$exit
      -- CP-element group 19: 	 branch_block_stmt_13736/assign_stmt_13743/RPIPE_e_cmd_pipe_13742_update_completed_
      -- CP-element group 19: 	 branch_block_stmt_13736/assign_stmt_13743/RPIPE_e_cmd_pipe_13742_Update/$exit
      -- CP-element group 19: 	 branch_block_stmt_13736/assign_stmt_13743/RPIPE_e_cmd_pipe_13742_Update/ca
      -- 
    ca_11172_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_e_cmd_pipe_13742_inst_ack_1, ack => e_block_daemon_CP_11105_elements(19)); -- 
    -- CP-element group 20:  join  fork  transition  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	4 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	5 
    -- CP-element group 20:  members (50) 
      -- CP-element group 20: 	 branch_block_stmt_13736/assign_stmt_13747_to_assign_stmt_13755/$entry
      -- CP-element group 20: 	 branch_block_stmt_13736/assign_stmt_13747_to_assign_stmt_13755/$exit
      -- CP-element group 20: 	 branch_block_stmt_13736/assign_stmt_13747_to_assign_stmt_13755/slice_13746_sample_start_
      -- CP-element group 20: 	 branch_block_stmt_13736/assign_stmt_13747_to_assign_stmt_13755/slice_13746_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_13736/assign_stmt_13747_to_assign_stmt_13755/slice_13746_update_start_
      -- CP-element group 20: 	 branch_block_stmt_13736/assign_stmt_13747_to_assign_stmt_13755/slice_13746_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_13736/assign_stmt_13747_to_assign_stmt_13755/R_e_init_cmd_13745_sample_start_
      -- CP-element group 20: 	 branch_block_stmt_13736/assign_stmt_13747_to_assign_stmt_13755/R_e_init_cmd_13745_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_13736/assign_stmt_13747_to_assign_stmt_13755/R_e_init_cmd_13745_update_start_
      -- CP-element group 20: 	 branch_block_stmt_13736/assign_stmt_13747_to_assign_stmt_13755/R_e_init_cmd_13745_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_13736/assign_stmt_13747_to_assign_stmt_13755/slice_13746_Sample/$entry
      -- CP-element group 20: 	 branch_block_stmt_13736/assign_stmt_13747_to_assign_stmt_13755/slice_13746_Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_13736/assign_stmt_13747_to_assign_stmt_13755/slice_13746_Sample/rr
      -- CP-element group 20: 	 branch_block_stmt_13736/assign_stmt_13747_to_assign_stmt_13755/slice_13746_Sample/ra
      -- CP-element group 20: 	 branch_block_stmt_13736/assign_stmt_13747_to_assign_stmt_13755/slice_13746_Update/$entry
      -- CP-element group 20: 	 branch_block_stmt_13736/assign_stmt_13747_to_assign_stmt_13755/slice_13746_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_13736/assign_stmt_13747_to_assign_stmt_13755/slice_13746_Update/cr
      -- CP-element group 20: 	 branch_block_stmt_13736/assign_stmt_13747_to_assign_stmt_13755/slice_13746_Update/ca
      -- CP-element group 20: 	 branch_block_stmt_13736/assign_stmt_13747_to_assign_stmt_13755/slice_13750_sample_start_
      -- CP-element group 20: 	 branch_block_stmt_13736/assign_stmt_13747_to_assign_stmt_13755/slice_13750_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_13736/assign_stmt_13747_to_assign_stmt_13755/slice_13750_update_start_
      -- CP-element group 20: 	 branch_block_stmt_13736/assign_stmt_13747_to_assign_stmt_13755/slice_13750_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_13736/assign_stmt_13747_to_assign_stmt_13755/R_e_init_cmd_13749_sample_start_
      -- CP-element group 20: 	 branch_block_stmt_13736/assign_stmt_13747_to_assign_stmt_13755/R_e_init_cmd_13749_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_13736/assign_stmt_13747_to_assign_stmt_13755/R_e_init_cmd_13749_update_start_
      -- CP-element group 20: 	 branch_block_stmt_13736/assign_stmt_13747_to_assign_stmt_13755/R_e_init_cmd_13749_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_13736/assign_stmt_13747_to_assign_stmt_13755/slice_13750_Sample/$entry
      -- CP-element group 20: 	 branch_block_stmt_13736/assign_stmt_13747_to_assign_stmt_13755/slice_13750_Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_13736/assign_stmt_13747_to_assign_stmt_13755/slice_13750_Sample/rr
      -- CP-element group 20: 	 branch_block_stmt_13736/assign_stmt_13747_to_assign_stmt_13755/slice_13750_Sample/ra
      -- CP-element group 20: 	 branch_block_stmt_13736/assign_stmt_13747_to_assign_stmt_13755/slice_13750_Update/$entry
      -- CP-element group 20: 	 branch_block_stmt_13736/assign_stmt_13747_to_assign_stmt_13755/slice_13750_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_13736/assign_stmt_13747_to_assign_stmt_13755/slice_13750_Update/cr
      -- CP-element group 20: 	 branch_block_stmt_13736/assign_stmt_13747_to_assign_stmt_13755/slice_13750_Update/ca
      -- CP-element group 20: 	 branch_block_stmt_13736/assign_stmt_13747_to_assign_stmt_13755/slice_13754_sample_start_
      -- CP-element group 20: 	 branch_block_stmt_13736/assign_stmt_13747_to_assign_stmt_13755/slice_13754_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_13736/assign_stmt_13747_to_assign_stmt_13755/slice_13754_update_start_
      -- CP-element group 20: 	 branch_block_stmt_13736/assign_stmt_13747_to_assign_stmt_13755/slice_13754_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_13736/assign_stmt_13747_to_assign_stmt_13755/R_e_init_cmd_13753_sample_start_
      -- CP-element group 20: 	 branch_block_stmt_13736/assign_stmt_13747_to_assign_stmt_13755/R_e_init_cmd_13753_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_13736/assign_stmt_13747_to_assign_stmt_13755/R_e_init_cmd_13753_update_start_
      -- CP-element group 20: 	 branch_block_stmt_13736/assign_stmt_13747_to_assign_stmt_13755/R_e_init_cmd_13753_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_13736/assign_stmt_13747_to_assign_stmt_13755/slice_13754_Sample/$entry
      -- CP-element group 20: 	 branch_block_stmt_13736/assign_stmt_13747_to_assign_stmt_13755/slice_13754_Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_13736/assign_stmt_13747_to_assign_stmt_13755/slice_13754_Sample/rr
      -- CP-element group 20: 	 branch_block_stmt_13736/assign_stmt_13747_to_assign_stmt_13755/slice_13754_Sample/ra
      -- CP-element group 20: 	 branch_block_stmt_13736/assign_stmt_13747_to_assign_stmt_13755/slice_13754_Update/$entry
      -- CP-element group 20: 	 branch_block_stmt_13736/assign_stmt_13747_to_assign_stmt_13755/slice_13754_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_13736/assign_stmt_13747_to_assign_stmt_13755/slice_13754_Update/cr
      -- CP-element group 20: 	 branch_block_stmt_13736/assign_stmt_13747_to_assign_stmt_13755/slice_13754_Update/ca
      -- 
    e_block_daemon_CP_11105_elements(20) <= e_block_daemon_CP_11105_elements(4);
    -- CP-element group 21:  transition  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	5 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_13736/if_stmt_13756_dead_link/$entry
      -- 
    e_block_daemon_CP_11105_elements(21) <= e_block_daemon_CP_11105_elements(5);
    -- CP-element group 22:  transition  output  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	5 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	23 
    -- CP-element group 22:  members (17) 
      -- CP-element group 22: 	 branch_block_stmt_13736/if_stmt_13756_eval_test/$entry
      -- CP-element group 22: 	 branch_block_stmt_13736/if_stmt_13756_eval_test/$exit
      -- CP-element group 22: 	 branch_block_stmt_13736/if_stmt_13756_eval_test/EQ_u1_u1_13759/$entry
      -- CP-element group 22: 	 branch_block_stmt_13736/if_stmt_13756_eval_test/EQ_u1_u1_13759/$exit
      -- CP-element group 22: 	 branch_block_stmt_13736/if_stmt_13756_eval_test/EQ_u1_u1_13759/EQ_u1_u1_13759_inputs/$entry
      -- CP-element group 22: 	 branch_block_stmt_13736/if_stmt_13756_eval_test/EQ_u1_u1_13759/EQ_u1_u1_13759_inputs/$exit
      -- CP-element group 22: 	 branch_block_stmt_13736/if_stmt_13756_eval_test/EQ_u1_u1_13759/SplitProtocol/$entry
      -- CP-element group 22: 	 branch_block_stmt_13736/if_stmt_13756_eval_test/EQ_u1_u1_13759/SplitProtocol/$exit
      -- CP-element group 22: 	 branch_block_stmt_13736/if_stmt_13756_eval_test/EQ_u1_u1_13759/SplitProtocol/Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_13736/if_stmt_13756_eval_test/EQ_u1_u1_13759/SplitProtocol/Sample/$exit
      -- CP-element group 22: 	 branch_block_stmt_13736/if_stmt_13756_eval_test/EQ_u1_u1_13759/SplitProtocol/Sample/rr
      -- CP-element group 22: 	 branch_block_stmt_13736/if_stmt_13756_eval_test/EQ_u1_u1_13759/SplitProtocol/Sample/ra
      -- CP-element group 22: 	 branch_block_stmt_13736/if_stmt_13756_eval_test/EQ_u1_u1_13759/SplitProtocol/Update/$entry
      -- CP-element group 22: 	 branch_block_stmt_13736/if_stmt_13756_eval_test/EQ_u1_u1_13759/SplitProtocol/Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_13736/if_stmt_13756_eval_test/EQ_u1_u1_13759/SplitProtocol/Update/cr
      -- CP-element group 22: 	 branch_block_stmt_13736/if_stmt_13756_eval_test/EQ_u1_u1_13759/SplitProtocol/Update/ca
      -- CP-element group 22: 	 branch_block_stmt_13736/if_stmt_13756_eval_test/branch_req
      -- 
    branch_req_11256_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_11256_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_block_daemon_CP_11105_elements(22), ack => if_stmt_13756_branch_req_0); -- 
    e_block_daemon_CP_11105_elements(22) <= e_block_daemon_CP_11105_elements(5);
    -- CP-element group 23:  branch  place  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	22 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	24 
    -- CP-element group 23: 	26 
    -- CP-element group 23:  members (1) 
      -- CP-element group 23: 	 branch_block_stmt_13736/EQ_u1_u1_13759_place
      -- 
    e_block_daemon_CP_11105_elements(23) <= e_block_daemon_CP_11105_elements(22);
    -- CP-element group 24:  transition  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	23 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24:  members (1) 
      -- CP-element group 24: 	 branch_block_stmt_13736/if_stmt_13756_if_link/$entry
      -- 
    e_block_daemon_CP_11105_elements(24) <= e_block_daemon_CP_11105_elements(23);
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	24 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	28 
    -- CP-element group 25:  members (2) 
      -- CP-element group 25: 	 branch_block_stmt_13736/if_stmt_13756_if_link/$exit
      -- CP-element group 25: 	 branch_block_stmt_13736/if_stmt_13756_if_link/if_choice_transition
      -- 
    if_choice_transition_11261_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_13756_branch_ack_1, ack => e_block_daemon_CP_11105_elements(25)); -- 
    -- CP-element group 26:  transition  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	23 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	27 
    -- CP-element group 26:  members (1) 
      -- CP-element group 26: 	 branch_block_stmt_13736/if_stmt_13756_else_link/$entry
      -- 
    e_block_daemon_CP_11105_elements(26) <= e_block_daemon_CP_11105_elements(23);
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	26 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	6 
    -- CP-element group 27:  members (2) 
      -- CP-element group 27: 	 branch_block_stmt_13736/if_stmt_13756_else_link/$exit
      -- CP-element group 27: 	 branch_block_stmt_13736/if_stmt_13756_else_link/else_choice_transition
      -- 
    else_choice_transition_11265_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_13756_branch_ack_0, ack => e_block_daemon_CP_11105_elements(27)); -- 
    -- CP-element group 28:  place  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	25 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	212 
    -- CP-element group 28:  members (1) 
      -- CP-element group 28: 	 branch_block_stmt_13736/NotGotCmd
      -- 
    e_block_daemon_CP_11105_elements(28) <= e_block_daemon_CP_11105_elements(25);
    -- CP-element group 29:  fork  transition  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	7 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29: 	31 
    -- CP-element group 29: 	33 
    -- CP-element group 29: 	35 
    -- CP-element group 29: 	37 
    -- CP-element group 29: 	39 
    -- CP-element group 29: 	41 
    -- CP-element group 29: 	43 
    -- CP-element group 29: 	45 
    -- CP-element group 29: 	47 
    -- CP-element group 29: 	49 
    -- CP-element group 29:  members (38) 
      -- CP-element group 29: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13811_Update/ccr
      -- CP-element group 29: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13816_update_start_
      -- CP-element group 29: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13816_Update/ccr
      -- CP-element group 29: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13816_Update/$entry
      -- CP-element group 29: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13821_update_start_
      -- CP-element group 29: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13811_Update/$entry
      -- CP-element group 29: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13821_Update/ccr
      -- CP-element group 29: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13821_Update/$entry
      -- CP-element group 29: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/$entry
      -- CP-element group 29: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13776_sample_start_
      -- CP-element group 29: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13776_update_start_
      -- CP-element group 29: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/R_K0_13772_sample_start_
      -- CP-element group 29: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/R_K0_13772_sample_completed_
      -- CP-element group 29: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/R_K0_13772_update_start_
      -- CP-element group 29: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/R_K0_13772_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13776_Sample/$entry
      -- CP-element group 29: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13776_Sample/crr
      -- CP-element group 29: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13776_Update/$entry
      -- CP-element group 29: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13776_Update/ccr
      -- CP-element group 29: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13781_update_start_
      -- CP-element group 29: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13781_Update/$entry
      -- CP-element group 29: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13781_Update/ccr
      -- CP-element group 29: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13786_update_start_
      -- CP-element group 29: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13786_Update/$entry
      -- CP-element group 29: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13786_Update/ccr
      -- CP-element group 29: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13791_update_start_
      -- CP-element group 29: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13791_Update/$entry
      -- CP-element group 29: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13791_Update/ccr
      -- CP-element group 29: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13796_update_start_
      -- CP-element group 29: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13796_Update/$entry
      -- CP-element group 29: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13796_Update/ccr
      -- CP-element group 29: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13801_update_start_
      -- CP-element group 29: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13801_Update/$entry
      -- CP-element group 29: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13801_Update/ccr
      -- CP-element group 29: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13806_update_start_
      -- CP-element group 29: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13806_Update/$entry
      -- CP-element group 29: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13806_Update/ccr
      -- CP-element group 29: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13811_update_start_
      -- 
    ccr_11286_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_11286_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_block_daemon_CP_11105_elements(29), ack => call_stmt_13776_call_req_1); -- 
    crr_11281_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_11281_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_block_daemon_CP_11105_elements(29), ack => call_stmt_13776_call_req_0); -- 
    ccr_11308_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_11308_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_block_daemon_CP_11105_elements(29), ack => call_stmt_13781_call_req_1); -- 
    ccr_11330_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_11330_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_block_daemon_CP_11105_elements(29), ack => call_stmt_13786_call_req_1); -- 
    ccr_11352_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_11352_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_block_daemon_CP_11105_elements(29), ack => call_stmt_13791_call_req_1); -- 
    ccr_11374_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_11374_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_block_daemon_CP_11105_elements(29), ack => call_stmt_13796_call_req_1); -- 
    ccr_11396_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_11396_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_block_daemon_CP_11105_elements(29), ack => call_stmt_13801_call_req_1); -- 
    ccr_11418_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_11418_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_block_daemon_CP_11105_elements(29), ack => call_stmt_13806_call_req_1); -- 
    ccr_11440_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_11440_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_block_daemon_CP_11105_elements(29), ack => call_stmt_13811_call_req_1); -- 
    ccr_11462_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_11462_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_block_daemon_CP_11105_elements(29), ack => call_stmt_13816_call_req_1); -- 
    ccr_11484_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_11484_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_block_daemon_CP_11105_elements(29), ack => call_stmt_13821_call_req_1); -- 
    e_block_daemon_CP_11105_elements(29) <= e_block_daemon_CP_11105_elements(7);
    -- CP-element group 30:  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13776_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13776_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13776_Sample/cra
      -- 
    cra_11282_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_13776_call_ack_0, ack => e_block_daemon_CP_11105_elements(30)); -- 
    -- CP-element group 31:  join  fork  transition  input  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	29 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31:  members (14) 
      -- CP-element group 31: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13776_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13776_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13776_Update/cca
      -- CP-element group 31: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13781_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/R_K1_13777_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/R_K1_13777_sample_completed_
      -- CP-element group 31: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/R_K1_13777_update_start_
      -- CP-element group 31: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/R_K1_13777_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/R_RConstant_2_13778_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/R_RConstant_2_13778_sample_completed_
      -- CP-element group 31: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/R_RConstant_2_13778_update_start_
      -- CP-element group 31: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/R_RConstant_2_13778_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13781_Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13781_Sample/crr
      -- 
    cca_11287_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_13776_call_ack_1, ack => e_block_daemon_CP_11105_elements(31)); -- 
    crr_11303_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_11303_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_block_daemon_CP_11105_elements(31), ack => call_stmt_13781_call_req_0); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13781_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13781_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13781_Sample/cra
      -- 
    cra_11304_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_13781_call_ack_0, ack => e_block_daemon_CP_11105_elements(32)); -- 
    -- CP-element group 33:  join  fork  transition  input  output  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	29 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (14) 
      -- CP-element group 33: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13781_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13781_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13781_Update/cca
      -- CP-element group 33: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13786_sample_start_
      -- CP-element group 33: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/R_K2_13782_sample_start_
      -- CP-element group 33: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/R_K2_13782_sample_completed_
      -- CP-element group 33: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/R_K2_13782_update_start_
      -- CP-element group 33: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/R_K2_13782_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/R_RConstant_3_13783_sample_start_
      -- CP-element group 33: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/R_RConstant_3_13783_sample_completed_
      -- CP-element group 33: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/R_RConstant_3_13783_update_start_
      -- CP-element group 33: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/R_RConstant_3_13783_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13786_Sample/$entry
      -- CP-element group 33: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13786_Sample/crr
      -- 
    cca_11309_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_13781_call_ack_1, ack => e_block_daemon_CP_11105_elements(33)); -- 
    crr_11325_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_11325_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_block_daemon_CP_11105_elements(33), ack => call_stmt_13786_call_req_0); -- 
    -- CP-element group 34:  transition  input  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13786_sample_completed_
      -- CP-element group 34: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13786_Sample/$exit
      -- CP-element group 34: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13786_Sample/cra
      -- 
    cra_11326_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_13786_call_ack_0, ack => e_block_daemon_CP_11105_elements(34)); -- 
    -- CP-element group 35:  join  fork  transition  input  output  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	29 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	36 
    -- CP-element group 35:  members (14) 
      -- CP-element group 35: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13786_update_completed_
      -- CP-element group 35: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13786_Update/$exit
      -- CP-element group 35: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13786_Update/cca
      -- CP-element group 35: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13791_sample_start_
      -- CP-element group 35: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/R_K3_13787_sample_start_
      -- CP-element group 35: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/R_K3_13787_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/R_K3_13787_update_start_
      -- CP-element group 35: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/R_K3_13787_update_completed_
      -- CP-element group 35: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/R_RConstant_4_13788_sample_start_
      -- CP-element group 35: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/R_RConstant_4_13788_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/R_RConstant_4_13788_update_start_
      -- CP-element group 35: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/R_RConstant_4_13788_update_completed_
      -- CP-element group 35: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13791_Sample/$entry
      -- CP-element group 35: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13791_Sample/crr
      -- 
    cca_11331_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_13786_call_ack_1, ack => e_block_daemon_CP_11105_elements(35)); -- 
    crr_11347_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_11347_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_block_daemon_CP_11105_elements(35), ack => call_stmt_13791_call_req_0); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	35 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13791_sample_completed_
      -- CP-element group 36: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13791_Sample/$exit
      -- CP-element group 36: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13791_Sample/cra
      -- 
    cra_11348_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_13791_call_ack_0, ack => e_block_daemon_CP_11105_elements(36)); -- 
    -- CP-element group 37:  join  fork  transition  input  output  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	29 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (14) 
      -- CP-element group 37: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13791_update_completed_
      -- CP-element group 37: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13791_Update/$exit
      -- CP-element group 37: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13791_Update/cca
      -- CP-element group 37: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13796_sample_start_
      -- CP-element group 37: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/R_K4_13792_sample_start_
      -- CP-element group 37: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/R_K4_13792_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/R_K4_13792_update_start_
      -- CP-element group 37: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/R_K4_13792_update_completed_
      -- CP-element group 37: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/R_RConstant_5_13793_sample_start_
      -- CP-element group 37: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/R_RConstant_5_13793_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/R_RConstant_5_13793_update_start_
      -- CP-element group 37: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/R_RConstant_5_13793_update_completed_
      -- CP-element group 37: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13796_Sample/$entry
      -- CP-element group 37: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13796_Sample/crr
      -- 
    cca_11353_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_13791_call_ack_1, ack => e_block_daemon_CP_11105_elements(37)); -- 
    crr_11369_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_11369_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_block_daemon_CP_11105_elements(37), ack => call_stmt_13796_call_req_0); -- 
    -- CP-element group 38:  transition  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13796_sample_completed_
      -- CP-element group 38: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13796_Sample/$exit
      -- CP-element group 38: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13796_Sample/cra
      -- 
    cra_11370_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_13796_call_ack_0, ack => e_block_daemon_CP_11105_elements(38)); -- 
    -- CP-element group 39:  join  fork  transition  input  output  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	29 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	40 
    -- CP-element group 39:  members (14) 
      -- CP-element group 39: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13796_update_completed_
      -- CP-element group 39: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13796_Update/$exit
      -- CP-element group 39: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13796_Update/cca
      -- CP-element group 39: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13801_sample_start_
      -- CP-element group 39: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/R_K5_13797_sample_start_
      -- CP-element group 39: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/R_K5_13797_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/R_K5_13797_update_start_
      -- CP-element group 39: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/R_K5_13797_update_completed_
      -- CP-element group 39: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/R_RConstant_6_13798_sample_start_
      -- CP-element group 39: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/R_RConstant_6_13798_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/R_RConstant_6_13798_update_start_
      -- CP-element group 39: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/R_RConstant_6_13798_update_completed_
      -- CP-element group 39: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13801_Sample/$entry
      -- CP-element group 39: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13801_Sample/crr
      -- 
    cca_11375_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_13796_call_ack_1, ack => e_block_daemon_CP_11105_elements(39)); -- 
    crr_11391_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_11391_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_block_daemon_CP_11105_elements(39), ack => call_stmt_13801_call_req_0); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	39 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13801_sample_completed_
      -- CP-element group 40: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13801_Sample/$exit
      -- CP-element group 40: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13801_Sample/cra
      -- 
    cra_11392_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_13801_call_ack_0, ack => e_block_daemon_CP_11105_elements(40)); -- 
    -- CP-element group 41:  join  fork  transition  input  output  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	29 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	42 
    -- CP-element group 41:  members (14) 
      -- CP-element group 41: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13801_update_completed_
      -- CP-element group 41: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13801_Update/$exit
      -- CP-element group 41: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13801_Update/cca
      -- CP-element group 41: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13806_sample_start_
      -- CP-element group 41: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/R_K6_13802_sample_start_
      -- CP-element group 41: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/R_K6_13802_sample_completed_
      -- CP-element group 41: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/R_K6_13802_update_start_
      -- CP-element group 41: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/R_K6_13802_update_completed_
      -- CP-element group 41: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/R_RConstant_7_13803_sample_start_
      -- CP-element group 41: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/R_RConstant_7_13803_sample_completed_
      -- CP-element group 41: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/R_RConstant_7_13803_update_start_
      -- CP-element group 41: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/R_RConstant_7_13803_update_completed_
      -- CP-element group 41: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13806_Sample/$entry
      -- CP-element group 41: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13806_Sample/crr
      -- 
    cca_11397_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_13801_call_ack_1, ack => e_block_daemon_CP_11105_elements(41)); -- 
    crr_11413_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_11413_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_block_daemon_CP_11105_elements(41), ack => call_stmt_13806_call_req_0); -- 
    -- CP-element group 42:  transition  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	41 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13806_sample_completed_
      -- CP-element group 42: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13806_Sample/$exit
      -- CP-element group 42: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13806_Sample/cra
      -- 
    cra_11414_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_13806_call_ack_0, ack => e_block_daemon_CP_11105_elements(42)); -- 
    -- CP-element group 43:  join  fork  transition  input  output  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	29 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	44 
    -- CP-element group 43:  members (14) 
      -- CP-element group 43: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13811_Sample/crr
      -- CP-element group 43: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13811_Sample/$entry
      -- CP-element group 43: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13806_update_completed_
      -- CP-element group 43: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13806_Update/$exit
      -- CP-element group 43: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13806_Update/cca
      -- CP-element group 43: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13811_sample_start_
      -- CP-element group 43: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/R_K7_13807_sample_start_
      -- CP-element group 43: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/R_K7_13807_sample_completed_
      -- CP-element group 43: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/R_K7_13807_update_start_
      -- CP-element group 43: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/R_K7_13807_update_completed_
      -- CP-element group 43: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/R_RConstant_8_13808_sample_start_
      -- CP-element group 43: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/R_RConstant_8_13808_sample_completed_
      -- CP-element group 43: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/R_RConstant_8_13808_update_start_
      -- CP-element group 43: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/R_RConstant_8_13808_update_completed_
      -- 
    cca_11419_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_13806_call_ack_1, ack => e_block_daemon_CP_11105_elements(43)); -- 
    crr_11435_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_11435_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_block_daemon_CP_11105_elements(43), ack => call_stmt_13811_call_req_0); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	43 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13811_Sample/cra
      -- CP-element group 44: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13811_Sample/$exit
      -- CP-element group 44: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13811_sample_completed_
      -- 
    cra_11436_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_13811_call_ack_0, ack => e_block_daemon_CP_11105_elements(44)); -- 
    -- CP-element group 45:  join  fork  transition  input  output  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	29 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45:  members (14) 
      -- CP-element group 45: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13811_Update/cca
      -- CP-element group 45: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/R_RConstant_9_13813_sample_completed_
      -- CP-element group 45: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/R_RConstant_9_13813_update_start_
      -- CP-element group 45: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13816_sample_start_
      -- CP-element group 45: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/R_K8_13812_sample_start_
      -- CP-element group 45: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/R_RConstant_9_13813_update_completed_
      -- CP-element group 45: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/R_K8_13812_sample_completed_
      -- CP-element group 45: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/R_K8_13812_update_start_
      -- CP-element group 45: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/R_K8_13812_update_completed_
      -- CP-element group 45: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13816_Sample/$entry
      -- CP-element group 45: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13816_Sample/crr
      -- CP-element group 45: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13811_Update/$exit
      -- CP-element group 45: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/R_RConstant_9_13813_sample_start_
      -- CP-element group 45: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13811_update_completed_
      -- 
    cca_11441_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_13811_call_ack_1, ack => e_block_daemon_CP_11105_elements(45)); -- 
    crr_11457_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_11457_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_block_daemon_CP_11105_elements(45), ack => call_stmt_13816_call_req_0); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13816_Sample/$exit
      -- CP-element group 46: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13816_Sample/cra
      -- CP-element group 46: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13816_sample_completed_
      -- 
    cra_11458_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_13816_call_ack_0, ack => e_block_daemon_CP_11105_elements(46)); -- 
    -- CP-element group 47:  join  fork  transition  input  output  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	29 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	48 
    -- CP-element group 47:  members (14) 
      -- CP-element group 47: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13816_Update/$exit
      -- CP-element group 47: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13816_update_completed_
      -- CP-element group 47: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13816_Update/cca
      -- CP-element group 47: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13821_sample_start_
      -- CP-element group 47: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/R_K9_13817_sample_start_
      -- CP-element group 47: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13821_Sample/crr
      -- CP-element group 47: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13821_Sample/$entry
      -- CP-element group 47: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/R_RConstant_10_13818_update_completed_
      -- CP-element group 47: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/R_RConstant_10_13818_update_start_
      -- CP-element group 47: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/R_RConstant_10_13818_sample_completed_
      -- CP-element group 47: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/R_RConstant_10_13818_sample_start_
      -- CP-element group 47: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/R_K9_13817_update_completed_
      -- CP-element group 47: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/R_K9_13817_update_start_
      -- CP-element group 47: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/R_K9_13817_sample_completed_
      -- 
    cca_11463_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_13816_call_ack_1, ack => e_block_daemon_CP_11105_elements(47)); -- 
    crr_11479_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_11479_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_block_daemon_CP_11105_elements(47), ack => call_stmt_13821_call_req_0); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	47 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13821_sample_completed_
      -- CP-element group 48: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13821_Sample/cra
      -- CP-element group 48: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13821_Sample/$exit
      -- 
    cra_11480_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_13821_call_ack_0, ack => e_block_daemon_CP_11105_elements(48)); -- 
    -- CP-element group 49:  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	29 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	8 
    -- CP-element group 49:  members (4) 
      -- CP-element group 49: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13821_Update/cca
      -- CP-element group 49: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13821_Update/$exit
      -- CP-element group 49: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/$exit
      -- CP-element group 49: 	 branch_block_stmt_13736/call_stmt_13776_to_call_stmt_13821/call_stmt_13821_update_completed_
      -- 
    cca_11485_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_13821_call_ack_1, ack => e_block_daemon_CP_11105_elements(49)); -- 
    -- CP-element group 50:  transition  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	9 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50:  members (1) 
      -- CP-element group 50: 	 branch_block_stmt_13736/do_while_stmt_13828/$entry
      -- 
    e_block_daemon_CP_11105_elements(50) <= e_block_daemon_CP_11105_elements(9);
    -- CP-element group 51:  place  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	57 
    -- CP-element group 51:  members (1) 
      -- CP-element group 51: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828__entry__
      -- 
    e_block_daemon_CP_11105_elements(51) <= e_block_daemon_CP_11105_elements(50);
    -- CP-element group 52:  merge  place  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	193 
    -- CP-element group 52:  members (1) 
      -- CP-element group 52: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828__exit__
      -- 
    -- Element group e_block_daemon_CP_11105_elements(52) is bound as output of CP function.
    -- CP-element group 53:  merge  place  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	56 
    -- CP-element group 53:  members (1) 
      -- CP-element group 53: 	 branch_block_stmt_13736/do_while_stmt_13828/loop_back
      -- 
    -- Element group e_block_daemon_CP_11105_elements(53) is bound as output of CP function.
    -- CP-element group 54:  branch  place  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	59 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	189 
    -- CP-element group 54: 	191 
    -- CP-element group 54:  members (1) 
      -- CP-element group 54: 	 branch_block_stmt_13736/do_while_stmt_13828/condition_done
      -- 
    e_block_daemon_CP_11105_elements(54) <= e_block_daemon_CP_11105_elements(59);
    -- CP-element group 55:  branch  place  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	249 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (1) 
      -- CP-element group 55: 	 branch_block_stmt_13736/do_while_stmt_13828/loop_body_done
      -- 
    e_block_daemon_CP_11105_elements(55) <= e_block_daemon_CP_11105_elements(249);
    -- CP-element group 56:  transition  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	53 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	64 
    -- CP-element group 56:  members (1) 
      -- CP-element group 56: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/back_edge_to_loop_body
      -- 
    e_block_daemon_CP_11105_elements(56) <= e_block_daemon_CP_11105_elements(53);
    -- CP-element group 57:  transition  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	51 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	66 
    -- CP-element group 57:  members (1) 
      -- CP-element group 57: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/first_time_through_loop_body
      -- 
    e_block_daemon_CP_11105_elements(57) <= e_block_daemon_CP_11105_elements(51);
    -- CP-element group 58:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	153 
    -- CP-element group 58: 	155 
    -- CP-element group 58: 	159 
    -- CP-element group 58: 	162 
    -- CP-element group 58: 	164 
    -- CP-element group 58: 	168 
    -- CP-element group 58: 	171 
    -- CP-element group 58: 	173 
    -- CP-element group 58: 	177 
    -- CP-element group 58: 	188 
    -- CP-element group 58: 	60 
    -- CP-element group 58: 	61 
    -- CP-element group 58: 	80 
    -- CP-element group 58: 	85 
    -- CP-element group 58: 	87 
    -- CP-element group 58: 	90 
    -- CP-element group 58: 	92 
    -- CP-element group 58: 	96 
    -- CP-element group 58: 	99 
    -- CP-element group 58: 	101 
    -- CP-element group 58: 	105 
    -- CP-element group 58: 	108 
    -- CP-element group 58: 	110 
    -- CP-element group 58: 	114 
    -- CP-element group 58: 	117 
    -- CP-element group 58: 	119 
    -- CP-element group 58: 	123 
    -- CP-element group 58: 	126 
    -- CP-element group 58: 	128 
    -- CP-element group 58: 	132 
    -- CP-element group 58: 	135 
    -- CP-element group 58: 	137 
    -- CP-element group 58: 	141 
    -- CP-element group 58: 	144 
    -- CP-element group 58: 	146 
    -- CP-element group 58: 	150 
    -- CP-element group 58:  members (28) 
      -- CP-element group 58: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_K1_13847_sample_completed_
      -- CP-element group 58: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_K1_13847_sample_start_
      -- CP-element group 58: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_K0_13840_sample_start_
      -- CP-element group 58: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/loop_body_start
      -- CP-element group 58: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/$entry
      -- CP-element group 58: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_K0_13840_sample_completed_
      -- CP-element group 58: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_K2_13855_sample_start_
      -- CP-element group 58: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_K2_13855_sample_completed_
      -- CP-element group 58: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_K3_13863_sample_start_
      -- CP-element group 58: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_K3_13863_sample_completed_
      -- CP-element group 58: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_K4_13871_sample_start_
      -- CP-element group 58: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_K4_13871_sample_completed_
      -- CP-element group 58: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_K5_13879_sample_start_
      -- CP-element group 58: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_K5_13879_sample_completed_
      -- CP-element group 58: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_K6_13887_sample_start_
      -- CP-element group 58: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_K6_13887_sample_completed_
      -- CP-element group 58: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_K7_13895_sample_start_
      -- CP-element group 58: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_K7_13895_sample_completed_
      -- CP-element group 58: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_K8_13903_sample_start_
      -- CP-element group 58: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_K8_13903_sample_completed_
      -- CP-element group 58: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_K9_13911_sample_start_
      -- CP-element group 58: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_K9_13911_sample_completed_
      -- CP-element group 58: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_K10_13919_sample_start_
      -- CP-element group 58: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_K10_13919_sample_completed_
      -- CP-element group 58: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_countB_13936_sample_start_
      -- CP-element group 58: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_countB_13936_sample_completed_
      -- CP-element group 58: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_countB_13936_update_start_
      -- CP-element group 58: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_countB_13936_update_completed_
      -- 
    -- Element group e_block_daemon_CP_11105_elements(58) is bound as output of CP function.
    -- CP-element group 59:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	188 
    -- CP-element group 59: 	61 
    -- CP-element group 59: 	62 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	54 
    -- CP-element group 59:  members (1) 
      -- CP-element group 59: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/condition_evaluated
      -- 
    condition_evaluated_11500_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_11500_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_block_daemon_CP_11105_elements(59), ack => do_while_stmt_13828_branch_req_0); -- 
    e_block_daemon_cp_element_group_59: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 2,1 => 2,2 => 2);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "e_block_daemon_cp_element_group_59"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= e_block_daemon_CP_11105_elements(188) & e_block_daemon_CP_11105_elements(61) & e_block_daemon_CP_11105_elements(62);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => e_block_daemon_CP_11105_elements(59), clk => clk, reset => reset); --
    end block;
    -- CP-element group 60:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	58 
    -- CP-element group 60: marked-predecessors 
    -- CP-element group 60: 	187 
    -- CP-element group 60: 	62 
    -- CP-element group 60: successors 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/phi_stmt_13830_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/phi_stmt_13830_sample_start__ps
      -- CP-element group 60: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/aggregated_phi_sample_req
      -- 
    e_block_daemon_cp_element_group_60: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 2,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 34) := "e_block_daemon_cp_element_group_60"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= e_block_daemon_CP_11105_elements(58) & e_block_daemon_CP_11105_elements(187) & e_block_daemon_CP_11105_elements(62);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => e_block_daemon_CP_11105_elements(60), clk => clk, reset => reset); --
    end block;
    -- CP-element group 61:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	58 
    -- CP-element group 61: marked-predecessors 
    -- CP-element group 61: 	186 
    -- CP-element group 61: 	63 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	59 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/aggregated_phi_update_req
      -- CP-element group 61: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/phi_stmt_13830_update_start_
      -- CP-element group 61: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/phi_stmt_13830_update_start__ps
      -- 
    e_block_daemon_cp_element_group_61: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 2,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "e_block_daemon_cp_element_group_61"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= e_block_daemon_CP_11105_elements(58) & e_block_daemon_CP_11105_elements(186) & e_block_daemon_CP_11105_elements(63);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => e_block_daemon_CP_11105_elements(61), clk => clk, reset => reset); --
    end block;
    -- CP-element group 62:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	185 
    -- CP-element group 62: 	59 
    -- CP-element group 62: marked-successors 
    -- CP-element group 62: 	60 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/phi_stmt_13830_sample_completed_
      -- CP-element group 62: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/aggregated_phi_sample_ack
      -- CP-element group 62: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/phi_stmt_13830_sample_completed__ps
      -- 
    -- Element group e_block_daemon_CP_11105_elements(62) is bound as output of CP function.
    -- CP-element group 63:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	184 
    -- CP-element group 63: marked-successors 
    -- CP-element group 63: 	61 
    -- CP-element group 63:  members (7) 
      -- CP-element group 63: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/aggregated_phi_update_ack
      -- CP-element group 63: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/phi_stmt_13830_update_completed_
      -- CP-element group 63: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/phi_stmt_13830_update_completed__ps
      -- CP-element group 63: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_count_var_13930_sample_start_
      -- CP-element group 63: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_count_var_13930_sample_completed_
      -- CP-element group 63: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_count_var_13930_update_start_
      -- CP-element group 63: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_count_var_13930_update_completed_
      -- 
    -- Element group e_block_daemon_CP_11105_elements(63) is bound as output of CP function.
    -- CP-element group 64:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	56 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (1) 
      -- CP-element group 64: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/phi_stmt_13830_loopback_trigger
      -- 
    e_block_daemon_CP_11105_elements(64) <= e_block_daemon_CP_11105_elements(56);
    -- CP-element group 65:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	70 
    -- CP-element group 65:  members (1) 
      -- CP-element group 65: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/phi_stmt_13830_loopback_sample_req
      -- 
    phi_stmt_13830_loopback_sample_req_11515_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_13830_loopback_sample_req_11515_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_block_daemon_CP_11105_elements(65), ack => phi_stmt_13830_req_1); -- 
    -- Element group e_block_daemon_CP_11105_elements(65) is bound as output of CP function.
    -- CP-element group 66:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	57 
    -- CP-element group 66: successors 
    -- CP-element group 66:  members (1) 
      -- CP-element group 66: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/phi_stmt_13830_entry_trigger
      -- 
    e_block_daemon_CP_11105_elements(66) <= e_block_daemon_CP_11105_elements(57);
    -- CP-element group 67:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	69 
    -- CP-element group 67:  members (1) 
      -- CP-element group 67: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/phi_stmt_13830_entry_sample_req
      -- 
    phi_stmt_13830_entry_sample_req_11517_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_13830_entry_sample_req_11517_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_block_daemon_CP_11105_elements(67), ack => phi_stmt_13830_req_0); -- 
    -- Element group e_block_daemon_CP_11105_elements(67) is bound as output of CP function.
    -- CP-element group 68:  transition  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: successors 
    -- CP-element group 68:  members (1) 
      -- CP-element group 68: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/phi_stmt_13830_merged_reqs
      -- 
    -- Element group e_block_daemon_CP_11105_elements(68) is bound as output of CP function.
    -- CP-element group 69:  transition  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	67 
    -- CP-element group 69: successors 
    -- CP-element group 69:  members (1) 
      -- CP-element group 69: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/phi_stmt_13830_entry_sample_req__merge_in
      -- 
    e_block_daemon_CP_11105_elements(69) <= e_block_daemon_CP_11105_elements(67);
    -- CP-element group 70:  transition  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	65 
    -- CP-element group 70: successors 
    -- CP-element group 70:  members (1) 
      -- CP-element group 70: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/phi_stmt_13830_loopback_sample_req__merge_in
      -- 
    e_block_daemon_CP_11105_elements(70) <= e_block_daemon_CP_11105_elements(65);
    -- CP-element group 71:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	249 
    -- CP-element group 71:  members (1) 
      -- CP-element group 71: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/phi_stmt_13830_phi_mux_ack
      -- 
    phi_stmt_13830_phi_mux_ack_11522_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_13830_ack_0, ack => e_block_daemon_CP_11105_elements(71)); -- 
    -- CP-element group 72:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: successors 
    -- CP-element group 72:  members (4) 
      -- CP-element group 72: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_ZERO_COUNT_13832_sample_completed_
      -- CP-element group 72: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_ZERO_COUNT_13832_sample_completed__ps
      -- CP-element group 72: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_ZERO_COUNT_13832_sample_start__ps
      -- CP-element group 72: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_ZERO_COUNT_13832_sample_start_
      -- 
    -- Element group e_block_daemon_CP_11105_elements(72) is bound as output of CP function.
    -- CP-element group 73:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	75 
    -- CP-element group 73:  members (2) 
      -- CP-element group 73: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_ZERO_COUNT_13832_update_start_
      -- CP-element group 73: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_ZERO_COUNT_13832_update_start__ps
      -- 
    -- Element group e_block_daemon_CP_11105_elements(73) is bound as output of CP function.
    -- CP-element group 74:  join  transition  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	75 
    -- CP-element group 74: successors 
    -- CP-element group 74:  members (1) 
      -- CP-element group 74: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_ZERO_COUNT_13832_update_completed__ps
      -- 
    e_block_daemon_CP_11105_elements(74) <= e_block_daemon_CP_11105_elements(75);
    -- CP-element group 75:  transition  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	73 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	74 
    -- CP-element group 75:  members (1) 
      -- CP-element group 75: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_ZERO_COUNT_13832_update_completed_
      -- 
    -- Element group e_block_daemon_CP_11105_elements(75) is a control-delay.
    cp_element_75_delay: control_delay_element  generic map(name => " 75_delay", delay_value => 1)  port map(req => e_block_daemon_CP_11105_elements(73), ack => e_block_daemon_CP_11105_elements(75), clk => clk, reset =>reset);
    -- CP-element group 76:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	78 
    -- CP-element group 76:  members (4) 
      -- CP-element group 76: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_n_count_var_13833_Sample/req
      -- CP-element group 76: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_n_count_var_13833_sample_start__ps
      -- CP-element group 76: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_n_count_var_13833_Sample/$entry
      -- CP-element group 76: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_n_count_var_13833_sample_start_
      -- 
    req_11543_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_11543_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_block_daemon_CP_11105_elements(76), ack => n_count_var_13933_13833_buf_req_0); -- 
    -- Element group e_block_daemon_CP_11105_elements(76) is bound as output of CP function.
    -- CP-element group 77:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	79 
    -- CP-element group 77:  members (4) 
      -- CP-element group 77: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_n_count_var_13833_update_start__ps
      -- CP-element group 77: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_n_count_var_13833_Update/req
      -- CP-element group 77: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_n_count_var_13833_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_n_count_var_13833_update_start_
      -- 
    req_11548_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_11548_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_block_daemon_CP_11105_elements(77), ack => n_count_var_13933_13833_buf_req_1); -- 
    -- Element group e_block_daemon_CP_11105_elements(77) is bound as output of CP function.
    -- CP-element group 78:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	76 
    -- CP-element group 78: successors 
    -- CP-element group 78:  members (4) 
      -- CP-element group 78: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_n_count_var_13833_Sample/$exit
      -- CP-element group 78: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_n_count_var_13833_sample_completed__ps
      -- CP-element group 78: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_n_count_var_13833_Sample/ack
      -- CP-element group 78: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_n_count_var_13833_sample_completed_
      -- 
    ack_11544_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_count_var_13933_13833_buf_ack_0, ack => e_block_daemon_CP_11105_elements(78)); -- 
    -- CP-element group 79:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	77 
    -- CP-element group 79: successors 
    -- CP-element group 79:  members (4) 
      -- CP-element group 79: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_n_count_var_13833_Update/ack
      -- CP-element group 79: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_n_count_var_13833_Update/$exit
      -- CP-element group 79: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_n_count_var_13833_update_completed_
      -- CP-element group 79: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_n_count_var_13833_update_completed__ps
      -- 
    ack_11549_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_count_var_13933_13833_buf_ack_1, ack => e_block_daemon_CP_11105_elements(79)); -- 
    -- CP-element group 80:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	58 
    -- CP-element group 80: marked-predecessors 
    -- CP-element group 80: 	82 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	82 
    -- CP-element group 80:  members (3) 
      -- CP-element group 80: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/RPIPE_e_in_buf_13836_Sample/rr
      -- CP-element group 80: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/RPIPE_e_in_buf_13836_Sample/$entry
      -- CP-element group 80: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/RPIPE_e_in_buf_13836_sample_start_
      -- 
    rr_11558_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11558_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_block_daemon_CP_11105_elements(80), ack => RPIPE_e_in_buf_13836_inst_req_0); -- 
    e_block_daemon_cp_element_group_80: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 2,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 34) := "e_block_daemon_cp_element_group_80"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= e_block_daemon_CP_11105_elements(58) & e_block_daemon_CP_11105_elements(82);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => e_block_daemon_CP_11105_elements(80), clk => clk, reset => reset); --
    end block;
    -- CP-element group 81:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	82 
    -- CP-element group 81: marked-predecessors 
    -- CP-element group 81: 	83 
    -- CP-element group 81: 	88 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	83 
    -- CP-element group 81:  members (3) 
      -- CP-element group 81: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/RPIPE_e_in_buf_13836_Update/cr
      -- CP-element group 81: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/RPIPE_e_in_buf_13836_Update/$entry
      -- CP-element group 81: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/RPIPE_e_in_buf_13836_update_start_
      -- 
    cr_11563_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11563_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_block_daemon_CP_11105_elements(81), ack => RPIPE_e_in_buf_13836_inst_req_1); -- 
    e_block_daemon_cp_element_group_81: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 2,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "e_block_daemon_cp_element_group_81"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= e_block_daemon_CP_11105_elements(82) & e_block_daemon_CP_11105_elements(83) & e_block_daemon_CP_11105_elements(88);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => e_block_daemon_CP_11105_elements(81), clk => clk, reset => reset); --
    end block;
    -- CP-element group 82:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	80 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	81 
    -- CP-element group 82: marked-successors 
    -- CP-element group 82: 	80 
    -- CP-element group 82:  members (3) 
      -- CP-element group 82: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/RPIPE_e_in_buf_13836_Sample/ra
      -- CP-element group 82: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/RPIPE_e_in_buf_13836_Sample/$exit
      -- CP-element group 82: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/RPIPE_e_in_buf_13836_sample_completed_
      -- 
    ra_11559_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_e_in_buf_13836_inst_ack_0, ack => e_block_daemon_CP_11105_elements(82)); -- 
    -- CP-element group 83:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	81 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	84 
    -- CP-element group 83: marked-successors 
    -- CP-element group 83: 	81 
    -- CP-element group 83:  members (7) 
      -- CP-element group 83: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/RPIPE_e_in_buf_13836_Update/$exit
      -- CP-element group 83: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_in128_13839_update_completed_
      -- CP-element group 83: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_in128_13839_update_start_
      -- CP-element group 83: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_in128_13839_sample_completed_
      -- CP-element group 83: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_in128_13839_sample_start_
      -- CP-element group 83: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/RPIPE_e_in_buf_13836_update_completed_
      -- CP-element group 83: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/RPIPE_e_in_buf_13836_Update/ca
      -- 
    ca_11564_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_e_in_buf_13836_inst_ack_1, ack => e_block_daemon_CP_11105_elements(83)); -- 
    -- CP-element group 84:  join  transition  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	83 
    -- CP-element group 84: 	85 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	86 
    -- CP-element group 84:  members (16) 
      -- CP-element group 84: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/XOR_u128_u128_13841_Update/ca
      -- CP-element group 84: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_round_S0_13844_update_completed_
      -- CP-element group 84: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_round_S0_13844_sample_start_
      -- CP-element group 84: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_round_S0_13844_update_start_
      -- CP-element group 84: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/XOR_u128_u128_13841_Update/cr
      -- CP-element group 84: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_round_S0_13844_sample_completed_
      -- CP-element group 84: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/XOR_u128_u128_13841_Update/$exit
      -- CP-element group 84: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/XOR_u128_u128_13841_Update/$entry
      -- CP-element group 84: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/XOR_u128_u128_13841_Sample/ra
      -- CP-element group 84: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/XOR_u128_u128_13841_Sample/rr
      -- CP-element group 84: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/XOR_u128_u128_13841_update_completed_
      -- CP-element group 84: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/XOR_u128_u128_13841_sample_completed_
      -- CP-element group 84: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/XOR_u128_u128_13841_Sample/$exit
      -- CP-element group 84: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/XOR_u128_u128_13841_Sample/$entry
      -- CP-element group 84: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/XOR_u128_u128_13841_update_start_
      -- CP-element group 84: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/XOR_u128_u128_13841_sample_start_
      -- 
    e_block_daemon_cp_element_group_84: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 2,1 => 2);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "e_block_daemon_cp_element_group_84"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= e_block_daemon_CP_11105_elements(83) & e_block_daemon_CP_11105_elements(85);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => e_block_daemon_CP_11105_elements(84), clk => clk, reset => reset); --
    end block;
    -- CP-element group 85:  join  transition  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	58 
    -- CP-element group 85: marked-predecessors 
    -- CP-element group 85: 	88 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	84 
    -- CP-element group 85:  members (2) 
      -- CP-element group 85: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_K0_13840_update_completed_
      -- CP-element group 85: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_K0_13840_update_start_
      -- 
    e_block_daemon_cp_element_group_85: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 2,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 34) := "e_block_daemon_cp_element_group_85"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= e_block_daemon_CP_11105_elements(58) & e_block_daemon_CP_11105_elements(88);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => e_block_daemon_CP_11105_elements(85), clk => clk, reset => reset); --
    end block;
    -- CP-element group 86:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	84 
    -- CP-element group 86: marked-predecessors 
    -- CP-element group 86: 	88 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	88 
    -- CP-element group 86:  members (3) 
      -- CP-element group 86: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13845_Sample/req
      -- CP-element group 86: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13845_sample_start_
      -- CP-element group 86: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13845_Sample/$entry
      -- 
    req_11598_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_11598_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_block_daemon_CP_11105_elements(86), ack => W_round_S0_13810_delayed_1_13843_inst_req_0); -- 
    e_block_daemon_cp_element_group_86: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 2,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 34) := "e_block_daemon_cp_element_group_86"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= e_block_daemon_CP_11105_elements(84) & e_block_daemon_CP_11105_elements(88);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => e_block_daemon_CP_11105_elements(86), clk => clk, reset => reset); --
    end block;
    -- CP-element group 87:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	58 
    -- CP-element group 87: marked-predecessors 
    -- CP-element group 87: 	89 
    -- CP-element group 87: 	97 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	89 
    -- CP-element group 87:  members (3) 
      -- CP-element group 87: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13845_Update/req
      -- CP-element group 87: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13845_Update/$entry
      -- CP-element group 87: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13845_update_start_
      -- 
    req_11603_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_11603_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_block_daemon_CP_11105_elements(87), ack => W_round_S0_13810_delayed_1_13843_inst_req_1); -- 
    e_block_daemon_cp_element_group_87: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 2,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "e_block_daemon_cp_element_group_87"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= e_block_daemon_CP_11105_elements(58) & e_block_daemon_CP_11105_elements(89) & e_block_daemon_CP_11105_elements(97);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => e_block_daemon_CP_11105_elements(87), clk => clk, reset => reset); --
    end block;
    -- CP-element group 88:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	86 
    -- CP-element group 88: successors 
    -- CP-element group 88: marked-successors 
    -- CP-element group 88: 	81 
    -- CP-element group 88: 	85 
    -- CP-element group 88: 	86 
    -- CP-element group 88:  members (3) 
      -- CP-element group 88: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13845_Sample/$exit
      -- CP-element group 88: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13845_Sample/ack
      -- CP-element group 88: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13845_sample_completed_
      -- 
    ack_11599_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_round_S0_13810_delayed_1_13843_inst_ack_0, ack => e_block_daemon_CP_11105_elements(88)); -- 
    -- CP-element group 89:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	87 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	95 
    -- CP-element group 89: marked-successors 
    -- CP-element group 89: 	87 
    -- CP-element group 89:  members (7) 
      -- CP-element group 89: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13845_Update/ack
      -- CP-element group 89: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13845_Update/$exit
      -- CP-element group 89: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13845_update_completed_
      -- CP-element group 89: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_round_S0_13810_delayed_1_13849_sample_start_
      -- CP-element group 89: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_round_S0_13810_delayed_1_13849_sample_completed_
      -- CP-element group 89: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_round_S0_13810_delayed_1_13849_update_start_
      -- CP-element group 89: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_round_S0_13810_delayed_1_13849_update_completed_
      -- 
    ack_11604_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_round_S0_13810_delayed_1_13843_inst_ack_1, ack => e_block_daemon_CP_11105_elements(89)); -- 
    -- CP-element group 90:  join  transition  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	58 
    -- CP-element group 90: marked-predecessors 
    -- CP-element group 90: 	93 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	91 
    -- CP-element group 90:  members (2) 
      -- CP-element group 90: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_K1_13847_update_start_
      -- CP-element group 90: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_K1_13847_update_completed_
      -- 
    e_block_daemon_cp_element_group_90: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 2,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 34) := "e_block_daemon_cp_element_group_90"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= e_block_daemon_CP_11105_elements(58) & e_block_daemon_CP_11105_elements(93);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => e_block_daemon_CP_11105_elements(90), clk => clk, reset => reset); --
    end block;
    -- CP-element group 91:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	90 
    -- CP-element group 91: marked-predecessors 
    -- CP-element group 91: 	93 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	93 
    -- CP-element group 91:  members (3) 
      -- CP-element group 91: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13848_sample_start_
      -- CP-element group 91: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13848_Sample/$entry
      -- CP-element group 91: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13848_Sample/req
      -- 
    req_11616_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_11616_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_block_daemon_CP_11105_elements(91), ack => W_K1_13811_delayed_1_13846_inst_req_0); -- 
    e_block_daemon_cp_element_group_91: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 2,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 34) := "e_block_daemon_cp_element_group_91"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= e_block_daemon_CP_11105_elements(90) & e_block_daemon_CP_11105_elements(93);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => e_block_daemon_CP_11105_elements(91), clk => clk, reset => reset); --
    end block;
    -- CP-element group 92:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	58 
    -- CP-element group 92: marked-predecessors 
    -- CP-element group 92: 	94 
    -- CP-element group 92: 	97 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	94 
    -- CP-element group 92:  members (3) 
      -- CP-element group 92: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13848_update_start_
      -- CP-element group 92: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13848_Update/$entry
      -- CP-element group 92: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13848_Update/req
      -- 
    req_11621_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_11621_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_block_daemon_CP_11105_elements(92), ack => W_K1_13811_delayed_1_13846_inst_req_1); -- 
    e_block_daemon_cp_element_group_92: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 2,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "e_block_daemon_cp_element_group_92"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= e_block_daemon_CP_11105_elements(58) & e_block_daemon_CP_11105_elements(94) & e_block_daemon_CP_11105_elements(97);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => e_block_daemon_CP_11105_elements(92), clk => clk, reset => reset); --
    end block;
    -- CP-element group 93:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	91 
    -- CP-element group 93: successors 
    -- CP-element group 93: marked-successors 
    -- CP-element group 93: 	90 
    -- CP-element group 93: 	91 
    -- CP-element group 93:  members (3) 
      -- CP-element group 93: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13848_sample_completed_
      -- CP-element group 93: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13848_Sample/$exit
      -- CP-element group 93: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13848_Sample/ack
      -- 
    ack_11617_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_K1_13811_delayed_1_13846_inst_ack_0, ack => e_block_daemon_CP_11105_elements(93)); -- 
    -- CP-element group 94:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	92 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	95 
    -- CP-element group 94: marked-successors 
    -- CP-element group 94: 	92 
    -- CP-element group 94:  members (7) 
      -- CP-element group 94: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13848_update_completed_
      -- CP-element group 94: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13848_Update/$exit
      -- CP-element group 94: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13848_Update/ack
      -- CP-element group 94: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_K1_13811_delayed_1_13850_sample_start_
      -- CP-element group 94: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_K1_13811_delayed_1_13850_sample_completed_
      -- CP-element group 94: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_K1_13811_delayed_1_13850_update_start_
      -- CP-element group 94: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_K1_13811_delayed_1_13850_update_completed_
      -- 
    ack_11622_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_K1_13811_delayed_1_13846_inst_ack_1, ack => e_block_daemon_CP_11105_elements(94)); -- 
    -- CP-element group 95:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	89 
    -- CP-element group 95: 	94 
    -- CP-element group 95: marked-predecessors 
    -- CP-element group 95: 	97 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	97 
    -- CP-element group 95:  members (3) 
      -- CP-element group 95: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13853_sample_start_
      -- CP-element group 95: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13853_Sample/$entry
      -- CP-element group 95: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13853_Sample/crr
      -- 
    crr_11638_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_11638_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_block_daemon_CP_11105_elements(95), ack => call_stmt_13853_call_req_0); -- 
    e_block_daemon_cp_element_group_95: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 2,1 => 2,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 34) := "e_block_daemon_cp_element_group_95"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= e_block_daemon_CP_11105_elements(89) & e_block_daemon_CP_11105_elements(94) & e_block_daemon_CP_11105_elements(97);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => e_block_daemon_CP_11105_elements(95), clk => clk, reset => reset); --
    end block;
    -- CP-element group 96:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	58 
    -- CP-element group 96: marked-predecessors 
    -- CP-element group 96: 	98 
    -- CP-element group 96: 	106 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	98 
    -- CP-element group 96:  members (3) 
      -- CP-element group 96: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13853_update_start_
      -- CP-element group 96: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13853_Update/$entry
      -- CP-element group 96: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13853_Update/ccr
      -- 
    ccr_11643_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_11643_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_block_daemon_CP_11105_elements(96), ack => call_stmt_13853_call_req_1); -- 
    e_block_daemon_cp_element_group_96: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 2,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "e_block_daemon_cp_element_group_96"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= e_block_daemon_CP_11105_elements(58) & e_block_daemon_CP_11105_elements(98) & e_block_daemon_CP_11105_elements(106);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => e_block_daemon_CP_11105_elements(96), clk => clk, reset => reset); --
    end block;
    -- CP-element group 97:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	95 
    -- CP-element group 97: successors 
    -- CP-element group 97: marked-successors 
    -- CP-element group 97: 	87 
    -- CP-element group 97: 	92 
    -- CP-element group 97: 	95 
    -- CP-element group 97:  members (3) 
      -- CP-element group 97: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13853_sample_completed_
      -- CP-element group 97: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13853_Sample/$exit
      -- CP-element group 97: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13853_Sample/cra
      -- 
    cra_11639_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_13853_call_ack_0, ack => e_block_daemon_CP_11105_elements(97)); -- 
    -- CP-element group 98:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	96 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	104 
    -- CP-element group 98: marked-successors 
    -- CP-element group 98: 	96 
    -- CP-element group 98:  members (7) 
      -- CP-element group 98: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13853_update_completed_
      -- CP-element group 98: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13853_Update/$exit
      -- CP-element group 98: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13853_Update/cca
      -- CP-element group 98: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_round_S1_13857_sample_start_
      -- CP-element group 98: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_round_S1_13857_sample_completed_
      -- CP-element group 98: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_round_S1_13857_update_start_
      -- CP-element group 98: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_round_S1_13857_update_completed_
      -- 
    cca_11644_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_13853_call_ack_1, ack => e_block_daemon_CP_11105_elements(98)); -- 
    -- CP-element group 99:  join  transition  bypass  pipeline-parent 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	58 
    -- CP-element group 99: marked-predecessors 
    -- CP-element group 99: 	102 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	100 
    -- CP-element group 99:  members (2) 
      -- CP-element group 99: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_K2_13855_update_start_
      -- CP-element group 99: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_K2_13855_update_completed_
      -- 
    e_block_daemon_cp_element_group_99: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 2,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 34) := "e_block_daemon_cp_element_group_99"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= e_block_daemon_CP_11105_elements(58) & e_block_daemon_CP_11105_elements(102);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => e_block_daemon_CP_11105_elements(99), clk => clk, reset => reset); --
    end block;
    -- CP-element group 100:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	99 
    -- CP-element group 100: marked-predecessors 
    -- CP-element group 100: 	102 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	102 
    -- CP-element group 100:  members (3) 
      -- CP-element group 100: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13856_sample_start_
      -- CP-element group 100: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13856_Sample/$entry
      -- CP-element group 100: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13856_Sample/req
      -- 
    req_11656_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_11656_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_block_daemon_CP_11105_elements(100), ack => W_K2_13816_delayed_2_13854_inst_req_0); -- 
    e_block_daemon_cp_element_group_100: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 2,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "e_block_daemon_cp_element_group_100"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= e_block_daemon_CP_11105_elements(99) & e_block_daemon_CP_11105_elements(102);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => e_block_daemon_CP_11105_elements(100), clk => clk, reset => reset); --
    end block;
    -- CP-element group 101:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	58 
    -- CP-element group 101: marked-predecessors 
    -- CP-element group 101: 	103 
    -- CP-element group 101: 	106 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	103 
    -- CP-element group 101:  members (3) 
      -- CP-element group 101: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13856_update_start_
      -- CP-element group 101: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13856_Update/$entry
      -- CP-element group 101: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13856_Update/req
      -- 
    req_11661_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_11661_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_block_daemon_CP_11105_elements(101), ack => W_K2_13816_delayed_2_13854_inst_req_1); -- 
    e_block_daemon_cp_element_group_101: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 2,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "e_block_daemon_cp_element_group_101"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= e_block_daemon_CP_11105_elements(58) & e_block_daemon_CP_11105_elements(103) & e_block_daemon_CP_11105_elements(106);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => e_block_daemon_CP_11105_elements(101), clk => clk, reset => reset); --
    end block;
    -- CP-element group 102:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	100 
    -- CP-element group 102: successors 
    -- CP-element group 102: marked-successors 
    -- CP-element group 102: 	99 
    -- CP-element group 102: 	100 
    -- CP-element group 102:  members (3) 
      -- CP-element group 102: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13856_sample_completed_
      -- CP-element group 102: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13856_Sample/$exit
      -- CP-element group 102: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13856_Sample/ack
      -- 
    ack_11657_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_K2_13816_delayed_2_13854_inst_ack_0, ack => e_block_daemon_CP_11105_elements(102)); -- 
    -- CP-element group 103:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	101 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	104 
    -- CP-element group 103: marked-successors 
    -- CP-element group 103: 	101 
    -- CP-element group 103:  members (7) 
      -- CP-element group 103: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13856_update_completed_
      -- CP-element group 103: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13856_Update/$exit
      -- CP-element group 103: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13856_Update/ack
      -- CP-element group 103: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_K2_13816_delayed_2_13858_sample_start_
      -- CP-element group 103: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_K2_13816_delayed_2_13858_sample_completed_
      -- CP-element group 103: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_K2_13816_delayed_2_13858_update_start_
      -- CP-element group 103: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_K2_13816_delayed_2_13858_update_completed_
      -- 
    ack_11662_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_K2_13816_delayed_2_13854_inst_ack_1, ack => e_block_daemon_CP_11105_elements(103)); -- 
    -- CP-element group 104:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	98 
    -- CP-element group 104: 	103 
    -- CP-element group 104: marked-predecessors 
    -- CP-element group 104: 	106 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	106 
    -- CP-element group 104:  members (3) 
      -- CP-element group 104: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13861_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13861_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13861_Sample/crr
      -- 
    crr_11678_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_11678_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_block_daemon_CP_11105_elements(104), ack => call_stmt_13861_call_req_0); -- 
    e_block_daemon_cp_element_group_104: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 2,1 => 2,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 35) := "e_block_daemon_cp_element_group_104"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= e_block_daemon_CP_11105_elements(98) & e_block_daemon_CP_11105_elements(103) & e_block_daemon_CP_11105_elements(106);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => e_block_daemon_CP_11105_elements(104), clk => clk, reset => reset); --
    end block;
    -- CP-element group 105:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	58 
    -- CP-element group 105: marked-predecessors 
    -- CP-element group 105: 	107 
    -- CP-element group 105: 	115 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	107 
    -- CP-element group 105:  members (3) 
      -- CP-element group 105: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13861_update_start_
      -- CP-element group 105: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13861_Update/$entry
      -- CP-element group 105: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13861_Update/ccr
      -- 
    ccr_11683_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_11683_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_block_daemon_CP_11105_elements(105), ack => call_stmt_13861_call_req_1); -- 
    e_block_daemon_cp_element_group_105: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 2,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "e_block_daemon_cp_element_group_105"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= e_block_daemon_CP_11105_elements(58) & e_block_daemon_CP_11105_elements(107) & e_block_daemon_CP_11105_elements(115);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => e_block_daemon_CP_11105_elements(105), clk => clk, reset => reset); --
    end block;
    -- CP-element group 106:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	104 
    -- CP-element group 106: successors 
    -- CP-element group 106: marked-successors 
    -- CP-element group 106: 	96 
    -- CP-element group 106: 	101 
    -- CP-element group 106: 	104 
    -- CP-element group 106:  members (3) 
      -- CP-element group 106: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13861_sample_completed_
      -- CP-element group 106: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13861_Sample/$exit
      -- CP-element group 106: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13861_Sample/cra
      -- 
    cra_11679_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_13861_call_ack_0, ack => e_block_daemon_CP_11105_elements(106)); -- 
    -- CP-element group 107:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	105 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	113 
    -- CP-element group 107: marked-successors 
    -- CP-element group 107: 	105 
    -- CP-element group 107:  members (7) 
      -- CP-element group 107: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13861_update_completed_
      -- CP-element group 107: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13861_Update/$exit
      -- CP-element group 107: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13861_Update/cca
      -- CP-element group 107: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_round_S2_13865_sample_start_
      -- CP-element group 107: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_round_S2_13865_sample_completed_
      -- CP-element group 107: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_round_S2_13865_update_start_
      -- CP-element group 107: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_round_S2_13865_update_completed_
      -- 
    cca_11684_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_13861_call_ack_1, ack => e_block_daemon_CP_11105_elements(107)); -- 
    -- CP-element group 108:  join  transition  bypass  pipeline-parent 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	58 
    -- CP-element group 108: marked-predecessors 
    -- CP-element group 108: 	111 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	109 
    -- CP-element group 108:  members (2) 
      -- CP-element group 108: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_K3_13863_update_start_
      -- CP-element group 108: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_K3_13863_update_completed_
      -- 
    e_block_daemon_cp_element_group_108: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 2,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "e_block_daemon_cp_element_group_108"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= e_block_daemon_CP_11105_elements(58) & e_block_daemon_CP_11105_elements(111);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => e_block_daemon_CP_11105_elements(108), clk => clk, reset => reset); --
    end block;
    -- CP-element group 109:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	108 
    -- CP-element group 109: marked-predecessors 
    -- CP-element group 109: 	111 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	111 
    -- CP-element group 109:  members (3) 
      -- CP-element group 109: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13864_Sample/$entry
      -- CP-element group 109: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13864_sample_start_
      -- CP-element group 109: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13864_Sample/req
      -- 
    req_11696_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_11696_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_block_daemon_CP_11105_elements(109), ack => W_K3_13821_delayed_3_13862_inst_req_0); -- 
    e_block_daemon_cp_element_group_109: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 2,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "e_block_daemon_cp_element_group_109"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= e_block_daemon_CP_11105_elements(108) & e_block_daemon_CP_11105_elements(111);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => e_block_daemon_CP_11105_elements(109), clk => clk, reset => reset); --
    end block;
    -- CP-element group 110:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	58 
    -- CP-element group 110: marked-predecessors 
    -- CP-element group 110: 	112 
    -- CP-element group 110: 	115 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	112 
    -- CP-element group 110:  members (3) 
      -- CP-element group 110: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13864_update_start_
      -- CP-element group 110: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13864_Update/$entry
      -- CP-element group 110: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13864_Update/req
      -- 
    req_11701_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_11701_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_block_daemon_CP_11105_elements(110), ack => W_K3_13821_delayed_3_13862_inst_req_1); -- 
    e_block_daemon_cp_element_group_110: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 2,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "e_block_daemon_cp_element_group_110"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= e_block_daemon_CP_11105_elements(58) & e_block_daemon_CP_11105_elements(112) & e_block_daemon_CP_11105_elements(115);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => e_block_daemon_CP_11105_elements(110), clk => clk, reset => reset); --
    end block;
    -- CP-element group 111:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	109 
    -- CP-element group 111: successors 
    -- CP-element group 111: marked-successors 
    -- CP-element group 111: 	108 
    -- CP-element group 111: 	109 
    -- CP-element group 111:  members (3) 
      -- CP-element group 111: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13864_sample_completed_
      -- CP-element group 111: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13864_Sample/$exit
      -- CP-element group 111: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13864_Sample/ack
      -- 
    ack_11697_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_K3_13821_delayed_3_13862_inst_ack_0, ack => e_block_daemon_CP_11105_elements(111)); -- 
    -- CP-element group 112:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	110 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	113 
    -- CP-element group 112: marked-successors 
    -- CP-element group 112: 	110 
    -- CP-element group 112:  members (7) 
      -- CP-element group 112: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13864_update_completed_
      -- CP-element group 112: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13864_Update/$exit
      -- CP-element group 112: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13864_Update/ack
      -- CP-element group 112: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_K3_13821_delayed_3_13866_sample_start_
      -- CP-element group 112: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_K3_13821_delayed_3_13866_sample_completed_
      -- CP-element group 112: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_K3_13821_delayed_3_13866_update_start_
      -- CP-element group 112: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_K3_13821_delayed_3_13866_update_completed_
      -- 
    ack_11702_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_K3_13821_delayed_3_13862_inst_ack_1, ack => e_block_daemon_CP_11105_elements(112)); -- 
    -- CP-element group 113:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	107 
    -- CP-element group 113: 	112 
    -- CP-element group 113: marked-predecessors 
    -- CP-element group 113: 	115 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	115 
    -- CP-element group 113:  members (3) 
      -- CP-element group 113: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13869_sample_start_
      -- CP-element group 113: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13869_Sample/$entry
      -- CP-element group 113: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13869_Sample/crr
      -- 
    crr_11718_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_11718_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_block_daemon_CP_11105_elements(113), ack => call_stmt_13869_call_req_0); -- 
    e_block_daemon_cp_element_group_113: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 2,1 => 2,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 35) := "e_block_daemon_cp_element_group_113"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= e_block_daemon_CP_11105_elements(107) & e_block_daemon_CP_11105_elements(112) & e_block_daemon_CP_11105_elements(115);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => e_block_daemon_CP_11105_elements(113), clk => clk, reset => reset); --
    end block;
    -- CP-element group 114:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	58 
    -- CP-element group 114: marked-predecessors 
    -- CP-element group 114: 	116 
    -- CP-element group 114: 	124 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	116 
    -- CP-element group 114:  members (3) 
      -- CP-element group 114: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13869_update_start_
      -- CP-element group 114: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13869_Update/$entry
      -- CP-element group 114: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13869_Update/ccr
      -- 
    ccr_11723_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_11723_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_block_daemon_CP_11105_elements(114), ack => call_stmt_13869_call_req_1); -- 
    e_block_daemon_cp_element_group_114: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 2,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "e_block_daemon_cp_element_group_114"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= e_block_daemon_CP_11105_elements(58) & e_block_daemon_CP_11105_elements(116) & e_block_daemon_CP_11105_elements(124);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => e_block_daemon_CP_11105_elements(114), clk => clk, reset => reset); --
    end block;
    -- CP-element group 115:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	113 
    -- CP-element group 115: successors 
    -- CP-element group 115: marked-successors 
    -- CP-element group 115: 	105 
    -- CP-element group 115: 	110 
    -- CP-element group 115: 	113 
    -- CP-element group 115:  members (3) 
      -- CP-element group 115: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13869_sample_completed_
      -- CP-element group 115: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13869_Sample/$exit
      -- CP-element group 115: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13869_Sample/cra
      -- 
    cra_11719_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_13869_call_ack_0, ack => e_block_daemon_CP_11105_elements(115)); -- 
    -- CP-element group 116:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	114 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	122 
    -- CP-element group 116: marked-successors 
    -- CP-element group 116: 	114 
    -- CP-element group 116:  members (7) 
      -- CP-element group 116: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13869_update_completed_
      -- CP-element group 116: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13869_Update/$exit
      -- CP-element group 116: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13869_Update/cca
      -- CP-element group 116: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_round_S3_13873_sample_start_
      -- CP-element group 116: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_round_S3_13873_sample_completed_
      -- CP-element group 116: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_round_S3_13873_update_start_
      -- CP-element group 116: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_round_S3_13873_update_completed_
      -- 
    cca_11724_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_13869_call_ack_1, ack => e_block_daemon_CP_11105_elements(116)); -- 
    -- CP-element group 117:  join  transition  bypass  pipeline-parent 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	58 
    -- CP-element group 117: marked-predecessors 
    -- CP-element group 117: 	120 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	118 
    -- CP-element group 117:  members (2) 
      -- CP-element group 117: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_K4_13871_update_start_
      -- CP-element group 117: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_K4_13871_update_completed_
      -- 
    e_block_daemon_cp_element_group_117: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 2,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "e_block_daemon_cp_element_group_117"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= e_block_daemon_CP_11105_elements(58) & e_block_daemon_CP_11105_elements(120);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => e_block_daemon_CP_11105_elements(117), clk => clk, reset => reset); --
    end block;
    -- CP-element group 118:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	117 
    -- CP-element group 118: marked-predecessors 
    -- CP-element group 118: 	120 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	120 
    -- CP-element group 118:  members (3) 
      -- CP-element group 118: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13872_sample_start_
      -- CP-element group 118: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13872_Sample/$entry
      -- CP-element group 118: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13872_Sample/req
      -- 
    req_11736_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_11736_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_block_daemon_CP_11105_elements(118), ack => W_K4_13826_delayed_4_13870_inst_req_0); -- 
    e_block_daemon_cp_element_group_118: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 2,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "e_block_daemon_cp_element_group_118"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= e_block_daemon_CP_11105_elements(117) & e_block_daemon_CP_11105_elements(120);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => e_block_daemon_CP_11105_elements(118), clk => clk, reset => reset); --
    end block;
    -- CP-element group 119:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	58 
    -- CP-element group 119: marked-predecessors 
    -- CP-element group 119: 	121 
    -- CP-element group 119: 	124 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	121 
    -- CP-element group 119:  members (3) 
      -- CP-element group 119: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13872_update_start_
      -- CP-element group 119: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13872_Update/$entry
      -- CP-element group 119: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13872_Update/req
      -- 
    req_11741_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_11741_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_block_daemon_CP_11105_elements(119), ack => W_K4_13826_delayed_4_13870_inst_req_1); -- 
    e_block_daemon_cp_element_group_119: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 2,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "e_block_daemon_cp_element_group_119"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= e_block_daemon_CP_11105_elements(58) & e_block_daemon_CP_11105_elements(121) & e_block_daemon_CP_11105_elements(124);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => e_block_daemon_CP_11105_elements(119), clk => clk, reset => reset); --
    end block;
    -- CP-element group 120:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	118 
    -- CP-element group 120: successors 
    -- CP-element group 120: marked-successors 
    -- CP-element group 120: 	117 
    -- CP-element group 120: 	118 
    -- CP-element group 120:  members (3) 
      -- CP-element group 120: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13872_sample_completed_
      -- CP-element group 120: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13872_Sample/$exit
      -- CP-element group 120: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13872_Sample/ack
      -- 
    ack_11737_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_K4_13826_delayed_4_13870_inst_ack_0, ack => e_block_daemon_CP_11105_elements(120)); -- 
    -- CP-element group 121:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	119 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	122 
    -- CP-element group 121: marked-successors 
    -- CP-element group 121: 	119 
    -- CP-element group 121:  members (7) 
      -- CP-element group 121: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13872_update_completed_
      -- CP-element group 121: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13872_Update/$exit
      -- CP-element group 121: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13872_Update/ack
      -- CP-element group 121: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_K4_13826_delayed_4_13874_sample_start_
      -- CP-element group 121: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_K4_13826_delayed_4_13874_sample_completed_
      -- CP-element group 121: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_K4_13826_delayed_4_13874_update_start_
      -- CP-element group 121: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_K4_13826_delayed_4_13874_update_completed_
      -- 
    ack_11742_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_K4_13826_delayed_4_13870_inst_ack_1, ack => e_block_daemon_CP_11105_elements(121)); -- 
    -- CP-element group 122:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	116 
    -- CP-element group 122: 	121 
    -- CP-element group 122: marked-predecessors 
    -- CP-element group 122: 	124 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	124 
    -- CP-element group 122:  members (3) 
      -- CP-element group 122: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13877_sample_start_
      -- CP-element group 122: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13877_Sample/$entry
      -- CP-element group 122: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13877_Sample/crr
      -- 
    crr_11758_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_11758_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_block_daemon_CP_11105_elements(122), ack => call_stmt_13877_call_req_0); -- 
    e_block_daemon_cp_element_group_122: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 2,1 => 2,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 35) := "e_block_daemon_cp_element_group_122"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= e_block_daemon_CP_11105_elements(116) & e_block_daemon_CP_11105_elements(121) & e_block_daemon_CP_11105_elements(124);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => e_block_daemon_CP_11105_elements(122), clk => clk, reset => reset); --
    end block;
    -- CP-element group 123:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	58 
    -- CP-element group 123: marked-predecessors 
    -- CP-element group 123: 	125 
    -- CP-element group 123: 	133 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	125 
    -- CP-element group 123:  members (3) 
      -- CP-element group 123: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13877_update_start_
      -- CP-element group 123: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13877_Update/$entry
      -- CP-element group 123: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13877_Update/ccr
      -- 
    ccr_11763_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_11763_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_block_daemon_CP_11105_elements(123), ack => call_stmt_13877_call_req_1); -- 
    e_block_daemon_cp_element_group_123: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 2,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "e_block_daemon_cp_element_group_123"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= e_block_daemon_CP_11105_elements(58) & e_block_daemon_CP_11105_elements(125) & e_block_daemon_CP_11105_elements(133);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => e_block_daemon_CP_11105_elements(123), clk => clk, reset => reset); --
    end block;
    -- CP-element group 124:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	122 
    -- CP-element group 124: successors 
    -- CP-element group 124: marked-successors 
    -- CP-element group 124: 	114 
    -- CP-element group 124: 	119 
    -- CP-element group 124: 	122 
    -- CP-element group 124:  members (3) 
      -- CP-element group 124: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13877_sample_completed_
      -- CP-element group 124: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13877_Sample/$exit
      -- CP-element group 124: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13877_Sample/cra
      -- 
    cra_11759_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_13877_call_ack_0, ack => e_block_daemon_CP_11105_elements(124)); -- 
    -- CP-element group 125:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	123 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	131 
    -- CP-element group 125: marked-successors 
    -- CP-element group 125: 	123 
    -- CP-element group 125:  members (7) 
      -- CP-element group 125: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13877_update_completed_
      -- CP-element group 125: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13877_Update/$exit
      -- CP-element group 125: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13877_Update/cca
      -- CP-element group 125: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_round_S4_13881_sample_start_
      -- CP-element group 125: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_round_S4_13881_sample_completed_
      -- CP-element group 125: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_round_S4_13881_update_start_
      -- CP-element group 125: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_round_S4_13881_update_completed_
      -- 
    cca_11764_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_13877_call_ack_1, ack => e_block_daemon_CP_11105_elements(125)); -- 
    -- CP-element group 126:  join  transition  bypass  pipeline-parent 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	58 
    -- CP-element group 126: marked-predecessors 
    -- CP-element group 126: 	129 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	127 
    -- CP-element group 126:  members (2) 
      -- CP-element group 126: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_K5_13879_update_start_
      -- CP-element group 126: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_K5_13879_update_completed_
      -- 
    e_block_daemon_cp_element_group_126: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 2,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "e_block_daemon_cp_element_group_126"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= e_block_daemon_CP_11105_elements(58) & e_block_daemon_CP_11105_elements(129);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => e_block_daemon_CP_11105_elements(126), clk => clk, reset => reset); --
    end block;
    -- CP-element group 127:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	126 
    -- CP-element group 127: marked-predecessors 
    -- CP-element group 127: 	129 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	129 
    -- CP-element group 127:  members (3) 
      -- CP-element group 127: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13880_sample_start_
      -- CP-element group 127: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13880_Sample/$entry
      -- CP-element group 127: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13880_Sample/req
      -- 
    req_11776_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_11776_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_block_daemon_CP_11105_elements(127), ack => W_K5_13831_delayed_5_13878_inst_req_0); -- 
    e_block_daemon_cp_element_group_127: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 2,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "e_block_daemon_cp_element_group_127"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= e_block_daemon_CP_11105_elements(126) & e_block_daemon_CP_11105_elements(129);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => e_block_daemon_CP_11105_elements(127), clk => clk, reset => reset); --
    end block;
    -- CP-element group 128:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	58 
    -- CP-element group 128: marked-predecessors 
    -- CP-element group 128: 	130 
    -- CP-element group 128: 	133 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	130 
    -- CP-element group 128:  members (3) 
      -- CP-element group 128: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13880_update_start_
      -- CP-element group 128: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13880_Update/$entry
      -- CP-element group 128: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13880_Update/req
      -- 
    req_11781_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_11781_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_block_daemon_CP_11105_elements(128), ack => W_K5_13831_delayed_5_13878_inst_req_1); -- 
    e_block_daemon_cp_element_group_128: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 2,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "e_block_daemon_cp_element_group_128"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= e_block_daemon_CP_11105_elements(58) & e_block_daemon_CP_11105_elements(130) & e_block_daemon_CP_11105_elements(133);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => e_block_daemon_CP_11105_elements(128), clk => clk, reset => reset); --
    end block;
    -- CP-element group 129:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	127 
    -- CP-element group 129: successors 
    -- CP-element group 129: marked-successors 
    -- CP-element group 129: 	126 
    -- CP-element group 129: 	127 
    -- CP-element group 129:  members (3) 
      -- CP-element group 129: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13880_sample_completed_
      -- CP-element group 129: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13880_Sample/$exit
      -- CP-element group 129: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13880_Sample/ack
      -- 
    ack_11777_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 129_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_K5_13831_delayed_5_13878_inst_ack_0, ack => e_block_daemon_CP_11105_elements(129)); -- 
    -- CP-element group 130:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	128 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	131 
    -- CP-element group 130: marked-successors 
    -- CP-element group 130: 	128 
    -- CP-element group 130:  members (7) 
      -- CP-element group 130: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13880_update_completed_
      -- CP-element group 130: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13880_Update/$exit
      -- CP-element group 130: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13880_Update/ack
      -- CP-element group 130: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_K5_13831_delayed_5_13882_sample_start_
      -- CP-element group 130: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_K5_13831_delayed_5_13882_sample_completed_
      -- CP-element group 130: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_K5_13831_delayed_5_13882_update_start_
      -- CP-element group 130: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_K5_13831_delayed_5_13882_update_completed_
      -- 
    ack_11782_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 130_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_K5_13831_delayed_5_13878_inst_ack_1, ack => e_block_daemon_CP_11105_elements(130)); -- 
    -- CP-element group 131:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	125 
    -- CP-element group 131: 	130 
    -- CP-element group 131: marked-predecessors 
    -- CP-element group 131: 	133 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	133 
    -- CP-element group 131:  members (3) 
      -- CP-element group 131: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13885_sample_start_
      -- CP-element group 131: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13885_Sample/$entry
      -- CP-element group 131: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13885_Sample/crr
      -- 
    crr_11798_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_11798_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_block_daemon_CP_11105_elements(131), ack => call_stmt_13885_call_req_0); -- 
    e_block_daemon_cp_element_group_131: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 2,1 => 2,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 35) := "e_block_daemon_cp_element_group_131"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= e_block_daemon_CP_11105_elements(125) & e_block_daemon_CP_11105_elements(130) & e_block_daemon_CP_11105_elements(133);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => e_block_daemon_CP_11105_elements(131), clk => clk, reset => reset); --
    end block;
    -- CP-element group 132:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	58 
    -- CP-element group 132: marked-predecessors 
    -- CP-element group 132: 	134 
    -- CP-element group 132: 	142 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	134 
    -- CP-element group 132:  members (3) 
      -- CP-element group 132: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13885_update_start_
      -- CP-element group 132: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13885_Update/$entry
      -- CP-element group 132: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13885_Update/ccr
      -- 
    ccr_11803_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_11803_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_block_daemon_CP_11105_elements(132), ack => call_stmt_13885_call_req_1); -- 
    e_block_daemon_cp_element_group_132: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 2,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "e_block_daemon_cp_element_group_132"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= e_block_daemon_CP_11105_elements(58) & e_block_daemon_CP_11105_elements(134) & e_block_daemon_CP_11105_elements(142);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => e_block_daemon_CP_11105_elements(132), clk => clk, reset => reset); --
    end block;
    -- CP-element group 133:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	131 
    -- CP-element group 133: successors 
    -- CP-element group 133: marked-successors 
    -- CP-element group 133: 	123 
    -- CP-element group 133: 	128 
    -- CP-element group 133: 	131 
    -- CP-element group 133:  members (3) 
      -- CP-element group 133: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13885_sample_completed_
      -- CP-element group 133: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13885_Sample/$exit
      -- CP-element group 133: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13885_Sample/cra
      -- 
    cra_11799_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_13885_call_ack_0, ack => e_block_daemon_CP_11105_elements(133)); -- 
    -- CP-element group 134:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	132 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	140 
    -- CP-element group 134: marked-successors 
    -- CP-element group 134: 	132 
    -- CP-element group 134:  members (7) 
      -- CP-element group 134: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13885_update_completed_
      -- CP-element group 134: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13885_Update/$exit
      -- CP-element group 134: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13885_Update/cca
      -- CP-element group 134: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_round_S5_13889_sample_start_
      -- CP-element group 134: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_round_S5_13889_sample_completed_
      -- CP-element group 134: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_round_S5_13889_update_start_
      -- CP-element group 134: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_round_S5_13889_update_completed_
      -- 
    cca_11804_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 134_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_13885_call_ack_1, ack => e_block_daemon_CP_11105_elements(134)); -- 
    -- CP-element group 135:  join  transition  bypass  pipeline-parent 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	58 
    -- CP-element group 135: marked-predecessors 
    -- CP-element group 135: 	138 
    -- CP-element group 135: successors 
    -- CP-element group 135: 	136 
    -- CP-element group 135:  members (2) 
      -- CP-element group 135: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_K6_13887_update_start_
      -- CP-element group 135: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_K6_13887_update_completed_
      -- 
    e_block_daemon_cp_element_group_135: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 2,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "e_block_daemon_cp_element_group_135"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= e_block_daemon_CP_11105_elements(58) & e_block_daemon_CP_11105_elements(138);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => e_block_daemon_CP_11105_elements(135), clk => clk, reset => reset); --
    end block;
    -- CP-element group 136:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	135 
    -- CP-element group 136: marked-predecessors 
    -- CP-element group 136: 	138 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	138 
    -- CP-element group 136:  members (3) 
      -- CP-element group 136: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13888_sample_start_
      -- CP-element group 136: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13888_Sample/$entry
      -- CP-element group 136: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13888_Sample/req
      -- 
    req_11816_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_11816_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_block_daemon_CP_11105_elements(136), ack => W_K6_13836_delayed_6_13886_inst_req_0); -- 
    e_block_daemon_cp_element_group_136: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 2,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "e_block_daemon_cp_element_group_136"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= e_block_daemon_CP_11105_elements(135) & e_block_daemon_CP_11105_elements(138);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => e_block_daemon_CP_11105_elements(136), clk => clk, reset => reset); --
    end block;
    -- CP-element group 137:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	58 
    -- CP-element group 137: marked-predecessors 
    -- CP-element group 137: 	139 
    -- CP-element group 137: 	142 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	139 
    -- CP-element group 137:  members (3) 
      -- CP-element group 137: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13888_update_start_
      -- CP-element group 137: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13888_Update/$entry
      -- CP-element group 137: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13888_Update/req
      -- 
    req_11821_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_11821_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_block_daemon_CP_11105_elements(137), ack => W_K6_13836_delayed_6_13886_inst_req_1); -- 
    e_block_daemon_cp_element_group_137: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 2,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "e_block_daemon_cp_element_group_137"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= e_block_daemon_CP_11105_elements(58) & e_block_daemon_CP_11105_elements(139) & e_block_daemon_CP_11105_elements(142);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => e_block_daemon_CP_11105_elements(137), clk => clk, reset => reset); --
    end block;
    -- CP-element group 138:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	136 
    -- CP-element group 138: successors 
    -- CP-element group 138: marked-successors 
    -- CP-element group 138: 	135 
    -- CP-element group 138: 	136 
    -- CP-element group 138:  members (3) 
      -- CP-element group 138: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13888_sample_completed_
      -- CP-element group 138: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13888_Sample/$exit
      -- CP-element group 138: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13888_Sample/ack
      -- 
    ack_11817_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 138_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_K6_13836_delayed_6_13886_inst_ack_0, ack => e_block_daemon_CP_11105_elements(138)); -- 
    -- CP-element group 139:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	137 
    -- CP-element group 139: successors 
    -- CP-element group 139: 	140 
    -- CP-element group 139: marked-successors 
    -- CP-element group 139: 	137 
    -- CP-element group 139:  members (7) 
      -- CP-element group 139: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13888_update_completed_
      -- CP-element group 139: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13888_Update/$exit
      -- CP-element group 139: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13888_Update/ack
      -- CP-element group 139: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_K6_13836_delayed_6_13890_sample_start_
      -- CP-element group 139: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_K6_13836_delayed_6_13890_sample_completed_
      -- CP-element group 139: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_K6_13836_delayed_6_13890_update_start_
      -- CP-element group 139: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_K6_13836_delayed_6_13890_update_completed_
      -- 
    ack_11822_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 139_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_K6_13836_delayed_6_13886_inst_ack_1, ack => e_block_daemon_CP_11105_elements(139)); -- 
    -- CP-element group 140:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	134 
    -- CP-element group 140: 	139 
    -- CP-element group 140: marked-predecessors 
    -- CP-element group 140: 	142 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	142 
    -- CP-element group 140:  members (3) 
      -- CP-element group 140: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13893_sample_start_
      -- CP-element group 140: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13893_Sample/$entry
      -- CP-element group 140: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13893_Sample/crr
      -- 
    crr_11838_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_11838_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_block_daemon_CP_11105_elements(140), ack => call_stmt_13893_call_req_0); -- 
    e_block_daemon_cp_element_group_140: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 2,1 => 2,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 35) := "e_block_daemon_cp_element_group_140"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= e_block_daemon_CP_11105_elements(134) & e_block_daemon_CP_11105_elements(139) & e_block_daemon_CP_11105_elements(142);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => e_block_daemon_CP_11105_elements(140), clk => clk, reset => reset); --
    end block;
    -- CP-element group 141:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	58 
    -- CP-element group 141: marked-predecessors 
    -- CP-element group 141: 	151 
    -- CP-element group 141: 	143 
    -- CP-element group 141: successors 
    -- CP-element group 141: 	143 
    -- CP-element group 141:  members (3) 
      -- CP-element group 141: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13893_update_start_
      -- CP-element group 141: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13893_Update/$entry
      -- CP-element group 141: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13893_Update/ccr
      -- 
    ccr_11843_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_11843_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_block_daemon_CP_11105_elements(141), ack => call_stmt_13893_call_req_1); -- 
    e_block_daemon_cp_element_group_141: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 2,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "e_block_daemon_cp_element_group_141"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= e_block_daemon_CP_11105_elements(58) & e_block_daemon_CP_11105_elements(151) & e_block_daemon_CP_11105_elements(143);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => e_block_daemon_CP_11105_elements(141), clk => clk, reset => reset); --
    end block;
    -- CP-element group 142:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	140 
    -- CP-element group 142: successors 
    -- CP-element group 142: marked-successors 
    -- CP-element group 142: 	132 
    -- CP-element group 142: 	137 
    -- CP-element group 142: 	140 
    -- CP-element group 142:  members (3) 
      -- CP-element group 142: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13893_sample_completed_
      -- CP-element group 142: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13893_Sample/$exit
      -- CP-element group 142: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13893_Sample/cra
      -- 
    cra_11839_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 142_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_13893_call_ack_0, ack => e_block_daemon_CP_11105_elements(142)); -- 
    -- CP-element group 143:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	141 
    -- CP-element group 143: successors 
    -- CP-element group 143: 	149 
    -- CP-element group 143: marked-successors 
    -- CP-element group 143: 	141 
    -- CP-element group 143:  members (7) 
      -- CP-element group 143: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13893_update_completed_
      -- CP-element group 143: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13893_Update/$exit
      -- CP-element group 143: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13893_Update/cca
      -- CP-element group 143: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_round_S6_13897_sample_start_
      -- CP-element group 143: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_round_S6_13897_sample_completed_
      -- CP-element group 143: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_round_S6_13897_update_start_
      -- CP-element group 143: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_round_S6_13897_update_completed_
      -- 
    cca_11844_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 143_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_13893_call_ack_1, ack => e_block_daemon_CP_11105_elements(143)); -- 
    -- CP-element group 144:  join  transition  bypass  pipeline-parent 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	58 
    -- CP-element group 144: marked-predecessors 
    -- CP-element group 144: 	147 
    -- CP-element group 144: successors 
    -- CP-element group 144: 	145 
    -- CP-element group 144:  members (2) 
      -- CP-element group 144: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_K7_13895_update_start_
      -- CP-element group 144: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_K7_13895_update_completed_
      -- 
    e_block_daemon_cp_element_group_144: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 2,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "e_block_daemon_cp_element_group_144"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= e_block_daemon_CP_11105_elements(58) & e_block_daemon_CP_11105_elements(147);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => e_block_daemon_CP_11105_elements(144), clk => clk, reset => reset); --
    end block;
    -- CP-element group 145:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	144 
    -- CP-element group 145: marked-predecessors 
    -- CP-element group 145: 	147 
    -- CP-element group 145: successors 
    -- CP-element group 145: 	147 
    -- CP-element group 145:  members (3) 
      -- CP-element group 145: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13896_sample_start_
      -- CP-element group 145: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13896_Sample/$entry
      -- CP-element group 145: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13896_Sample/req
      -- 
    req_11856_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_11856_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_block_daemon_CP_11105_elements(145), ack => W_K7_13841_delayed_7_13894_inst_req_0); -- 
    e_block_daemon_cp_element_group_145: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 2,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "e_block_daemon_cp_element_group_145"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= e_block_daemon_CP_11105_elements(144) & e_block_daemon_CP_11105_elements(147);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => e_block_daemon_CP_11105_elements(145), clk => clk, reset => reset); --
    end block;
    -- CP-element group 146:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	58 
    -- CP-element group 146: marked-predecessors 
    -- CP-element group 146: 	151 
    -- CP-element group 146: 	148 
    -- CP-element group 146: successors 
    -- CP-element group 146: 	148 
    -- CP-element group 146:  members (3) 
      -- CP-element group 146: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13896_update_start_
      -- CP-element group 146: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13896_Update/$entry
      -- CP-element group 146: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13896_Update/req
      -- 
    req_11861_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_11861_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_block_daemon_CP_11105_elements(146), ack => W_K7_13841_delayed_7_13894_inst_req_1); -- 
    e_block_daemon_cp_element_group_146: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 2,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "e_block_daemon_cp_element_group_146"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= e_block_daemon_CP_11105_elements(58) & e_block_daemon_CP_11105_elements(151) & e_block_daemon_CP_11105_elements(148);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => e_block_daemon_CP_11105_elements(146), clk => clk, reset => reset); --
    end block;
    -- CP-element group 147:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	145 
    -- CP-element group 147: successors 
    -- CP-element group 147: marked-successors 
    -- CP-element group 147: 	144 
    -- CP-element group 147: 	145 
    -- CP-element group 147:  members (3) 
      -- CP-element group 147: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13896_sample_completed_
      -- CP-element group 147: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13896_Sample/$exit
      -- CP-element group 147: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13896_Sample/ack
      -- 
    ack_11857_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 147_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_K7_13841_delayed_7_13894_inst_ack_0, ack => e_block_daemon_CP_11105_elements(147)); -- 
    -- CP-element group 148:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	146 
    -- CP-element group 148: successors 
    -- CP-element group 148: 	149 
    -- CP-element group 148: marked-successors 
    -- CP-element group 148: 	146 
    -- CP-element group 148:  members (7) 
      -- CP-element group 148: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13896_update_completed_
      -- CP-element group 148: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13896_Update/$exit
      -- CP-element group 148: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13896_Update/ack
      -- CP-element group 148: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_K7_13841_delayed_7_13898_sample_start_
      -- CP-element group 148: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_K7_13841_delayed_7_13898_sample_completed_
      -- CP-element group 148: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_K7_13841_delayed_7_13898_update_start_
      -- CP-element group 148: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_K7_13841_delayed_7_13898_update_completed_
      -- 
    ack_11862_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 148_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_K7_13841_delayed_7_13894_inst_ack_1, ack => e_block_daemon_CP_11105_elements(148)); -- 
    -- CP-element group 149:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	143 
    -- CP-element group 149: 	148 
    -- CP-element group 149: marked-predecessors 
    -- CP-element group 149: 	151 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	151 
    -- CP-element group 149:  members (3) 
      -- CP-element group 149: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13901_sample_start_
      -- CP-element group 149: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13901_Sample/$entry
      -- CP-element group 149: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13901_Sample/crr
      -- 
    crr_11878_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_11878_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_block_daemon_CP_11105_elements(149), ack => call_stmt_13901_call_req_0); -- 
    e_block_daemon_cp_element_group_149: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 2,1 => 2,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 35) := "e_block_daemon_cp_element_group_149"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= e_block_daemon_CP_11105_elements(143) & e_block_daemon_CP_11105_elements(148) & e_block_daemon_CP_11105_elements(151);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => e_block_daemon_CP_11105_elements(149), clk => clk, reset => reset); --
    end block;
    -- CP-element group 150:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	58 
    -- CP-element group 150: marked-predecessors 
    -- CP-element group 150: 	152 
    -- CP-element group 150: 	160 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	152 
    -- CP-element group 150:  members (3) 
      -- CP-element group 150: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13901_update_start_
      -- CP-element group 150: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13901_Update/$entry
      -- CP-element group 150: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13901_Update/ccr
      -- 
    ccr_11883_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_11883_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_block_daemon_CP_11105_elements(150), ack => call_stmt_13901_call_req_1); -- 
    e_block_daemon_cp_element_group_150: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 2,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "e_block_daemon_cp_element_group_150"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= e_block_daemon_CP_11105_elements(58) & e_block_daemon_CP_11105_elements(152) & e_block_daemon_CP_11105_elements(160);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => e_block_daemon_CP_11105_elements(150), clk => clk, reset => reset); --
    end block;
    -- CP-element group 151:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	149 
    -- CP-element group 151: successors 
    -- CP-element group 151: marked-successors 
    -- CP-element group 151: 	141 
    -- CP-element group 151: 	146 
    -- CP-element group 151: 	149 
    -- CP-element group 151:  members (3) 
      -- CP-element group 151: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13901_sample_completed_
      -- CP-element group 151: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13901_Sample/$exit
      -- CP-element group 151: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13901_Sample/cra
      -- 
    cra_11879_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 151_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_13901_call_ack_0, ack => e_block_daemon_CP_11105_elements(151)); -- 
    -- CP-element group 152:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	150 
    -- CP-element group 152: successors 
    -- CP-element group 152: 	158 
    -- CP-element group 152: marked-successors 
    -- CP-element group 152: 	150 
    -- CP-element group 152:  members (7) 
      -- CP-element group 152: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_round_S7_13905_update_start_
      -- CP-element group 152: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_round_S7_13905_update_completed_
      -- CP-element group 152: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13901_update_completed_
      -- CP-element group 152: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13901_Update/$exit
      -- CP-element group 152: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13901_Update/cca
      -- CP-element group 152: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_round_S7_13905_sample_start_
      -- CP-element group 152: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_round_S7_13905_sample_completed_
      -- 
    cca_11884_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_13901_call_ack_1, ack => e_block_daemon_CP_11105_elements(152)); -- 
    -- CP-element group 153:  join  transition  bypass  pipeline-parent 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	58 
    -- CP-element group 153: marked-predecessors 
    -- CP-element group 153: 	156 
    -- CP-element group 153: successors 
    -- CP-element group 153: 	154 
    -- CP-element group 153:  members (2) 
      -- CP-element group 153: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_K8_13903_update_start_
      -- CP-element group 153: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_K8_13903_update_completed_
      -- 
    e_block_daemon_cp_element_group_153: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 2,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "e_block_daemon_cp_element_group_153"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= e_block_daemon_CP_11105_elements(58) & e_block_daemon_CP_11105_elements(156);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => e_block_daemon_CP_11105_elements(153), clk => clk, reset => reset); --
    end block;
    -- CP-element group 154:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	153 
    -- CP-element group 154: marked-predecessors 
    -- CP-element group 154: 	156 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	156 
    -- CP-element group 154:  members (3) 
      -- CP-element group 154: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13904_sample_start_
      -- CP-element group 154: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13904_Sample/$entry
      -- CP-element group 154: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13904_Sample/req
      -- 
    req_11896_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_11896_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_block_daemon_CP_11105_elements(154), ack => W_K8_13846_delayed_8_13902_inst_req_0); -- 
    e_block_daemon_cp_element_group_154: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 2,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "e_block_daemon_cp_element_group_154"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= e_block_daemon_CP_11105_elements(153) & e_block_daemon_CP_11105_elements(156);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => e_block_daemon_CP_11105_elements(154), clk => clk, reset => reset); --
    end block;
    -- CP-element group 155:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	58 
    -- CP-element group 155: marked-predecessors 
    -- CP-element group 155: 	157 
    -- CP-element group 155: 	160 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	157 
    -- CP-element group 155:  members (3) 
      -- CP-element group 155: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13904_update_start_
      -- CP-element group 155: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13904_Update/$entry
      -- CP-element group 155: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13904_Update/req
      -- 
    req_11901_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_11901_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_block_daemon_CP_11105_elements(155), ack => W_K8_13846_delayed_8_13902_inst_req_1); -- 
    e_block_daemon_cp_element_group_155: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 2,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "e_block_daemon_cp_element_group_155"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= e_block_daemon_CP_11105_elements(58) & e_block_daemon_CP_11105_elements(157) & e_block_daemon_CP_11105_elements(160);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => e_block_daemon_CP_11105_elements(155), clk => clk, reset => reset); --
    end block;
    -- CP-element group 156:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	154 
    -- CP-element group 156: successors 
    -- CP-element group 156: marked-successors 
    -- CP-element group 156: 	153 
    -- CP-element group 156: 	154 
    -- CP-element group 156:  members (3) 
      -- CP-element group 156: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13904_sample_completed_
      -- CP-element group 156: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13904_Sample/$exit
      -- CP-element group 156: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13904_Sample/ack
      -- 
    ack_11897_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 156_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_K8_13846_delayed_8_13902_inst_ack_0, ack => e_block_daemon_CP_11105_elements(156)); -- 
    -- CP-element group 157:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	155 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	158 
    -- CP-element group 157: marked-successors 
    -- CP-element group 157: 	155 
    -- CP-element group 157:  members (7) 
      -- CP-element group 157: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13904_update_completed_
      -- CP-element group 157: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13904_Update/$exit
      -- CP-element group 157: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13904_Update/ack
      -- CP-element group 157: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_K8_13846_delayed_8_13906_sample_start_
      -- CP-element group 157: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_K8_13846_delayed_8_13906_sample_completed_
      -- CP-element group 157: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_K8_13846_delayed_8_13906_update_start_
      -- CP-element group 157: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_K8_13846_delayed_8_13906_update_completed_
      -- 
    ack_11902_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 157_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_K8_13846_delayed_8_13902_inst_ack_1, ack => e_block_daemon_CP_11105_elements(157)); -- 
    -- CP-element group 158:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	152 
    -- CP-element group 158: 	157 
    -- CP-element group 158: marked-predecessors 
    -- CP-element group 158: 	160 
    -- CP-element group 158: successors 
    -- CP-element group 158: 	160 
    -- CP-element group 158:  members (3) 
      -- CP-element group 158: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13909_sample_start_
      -- CP-element group 158: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13909_Sample/$entry
      -- CP-element group 158: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13909_Sample/crr
      -- 
    crr_11918_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_11918_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_block_daemon_CP_11105_elements(158), ack => call_stmt_13909_call_req_0); -- 
    e_block_daemon_cp_element_group_158: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 2,1 => 2,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 35) := "e_block_daemon_cp_element_group_158"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= e_block_daemon_CP_11105_elements(152) & e_block_daemon_CP_11105_elements(157) & e_block_daemon_CP_11105_elements(160);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => e_block_daemon_CP_11105_elements(158), clk => clk, reset => reset); --
    end block;
    -- CP-element group 159:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	58 
    -- CP-element group 159: marked-predecessors 
    -- CP-element group 159: 	161 
    -- CP-element group 159: 	169 
    -- CP-element group 159: successors 
    -- CP-element group 159: 	161 
    -- CP-element group 159:  members (3) 
      -- CP-element group 159: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13909_update_start_
      -- CP-element group 159: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13909_Update/$entry
      -- CP-element group 159: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13909_Update/ccr
      -- 
    ccr_11923_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_11923_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_block_daemon_CP_11105_elements(159), ack => call_stmt_13909_call_req_1); -- 
    e_block_daemon_cp_element_group_159: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 2,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "e_block_daemon_cp_element_group_159"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= e_block_daemon_CP_11105_elements(58) & e_block_daemon_CP_11105_elements(161) & e_block_daemon_CP_11105_elements(169);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => e_block_daemon_CP_11105_elements(159), clk => clk, reset => reset); --
    end block;
    -- CP-element group 160:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	158 
    -- CP-element group 160: successors 
    -- CP-element group 160: marked-successors 
    -- CP-element group 160: 	155 
    -- CP-element group 160: 	158 
    -- CP-element group 160: 	150 
    -- CP-element group 160:  members (3) 
      -- CP-element group 160: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13909_sample_completed_
      -- CP-element group 160: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13909_Sample/$exit
      -- CP-element group 160: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13909_Sample/cra
      -- 
    cra_11919_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 160_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_13909_call_ack_0, ack => e_block_daemon_CP_11105_elements(160)); -- 
    -- CP-element group 161:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	159 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	167 
    -- CP-element group 161: marked-successors 
    -- CP-element group 161: 	159 
    -- CP-element group 161:  members (7) 
      -- CP-element group 161: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13909_update_completed_
      -- CP-element group 161: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13909_Update/$exit
      -- CP-element group 161: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13909_Update/cca
      -- CP-element group 161: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_round_S8_13913_sample_start_
      -- CP-element group 161: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_round_S8_13913_sample_completed_
      -- CP-element group 161: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_round_S8_13913_update_start_
      -- CP-element group 161: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_round_S8_13913_update_completed_
      -- 
    cca_11924_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 161_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_13909_call_ack_1, ack => e_block_daemon_CP_11105_elements(161)); -- 
    -- CP-element group 162:  join  transition  bypass  pipeline-parent 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	58 
    -- CP-element group 162: marked-predecessors 
    -- CP-element group 162: 	165 
    -- CP-element group 162: successors 
    -- CP-element group 162: 	163 
    -- CP-element group 162:  members (2) 
      -- CP-element group 162: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_K9_13911_update_start_
      -- CP-element group 162: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_K9_13911_update_completed_
      -- 
    e_block_daemon_cp_element_group_162: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 2,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "e_block_daemon_cp_element_group_162"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= e_block_daemon_CP_11105_elements(58) & e_block_daemon_CP_11105_elements(165);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => e_block_daemon_CP_11105_elements(162), clk => clk, reset => reset); --
    end block;
    -- CP-element group 163:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	162 
    -- CP-element group 163: marked-predecessors 
    -- CP-element group 163: 	165 
    -- CP-element group 163: successors 
    -- CP-element group 163: 	165 
    -- CP-element group 163:  members (3) 
      -- CP-element group 163: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13912_sample_start_
      -- CP-element group 163: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13912_Sample/$entry
      -- CP-element group 163: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13912_Sample/req
      -- 
    req_11936_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_11936_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_block_daemon_CP_11105_elements(163), ack => W_K9_13851_delayed_9_13910_inst_req_0); -- 
    e_block_daemon_cp_element_group_163: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 2,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "e_block_daemon_cp_element_group_163"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= e_block_daemon_CP_11105_elements(162) & e_block_daemon_CP_11105_elements(165);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => e_block_daemon_CP_11105_elements(163), clk => clk, reset => reset); --
    end block;
    -- CP-element group 164:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: 	58 
    -- CP-element group 164: marked-predecessors 
    -- CP-element group 164: 	166 
    -- CP-element group 164: 	169 
    -- CP-element group 164: successors 
    -- CP-element group 164: 	166 
    -- CP-element group 164:  members (3) 
      -- CP-element group 164: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13912_update_start_
      -- CP-element group 164: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13912_Update/$entry
      -- CP-element group 164: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13912_Update/req
      -- 
    req_11941_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_11941_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_block_daemon_CP_11105_elements(164), ack => W_K9_13851_delayed_9_13910_inst_req_1); -- 
    e_block_daemon_cp_element_group_164: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 2,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "e_block_daemon_cp_element_group_164"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= e_block_daemon_CP_11105_elements(58) & e_block_daemon_CP_11105_elements(166) & e_block_daemon_CP_11105_elements(169);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => e_block_daemon_CP_11105_elements(164), clk => clk, reset => reset); --
    end block;
    -- CP-element group 165:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	163 
    -- CP-element group 165: successors 
    -- CP-element group 165: marked-successors 
    -- CP-element group 165: 	162 
    -- CP-element group 165: 	163 
    -- CP-element group 165:  members (3) 
      -- CP-element group 165: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13912_sample_completed_
      -- CP-element group 165: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13912_Sample/$exit
      -- CP-element group 165: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13912_Sample/ack
      -- 
    ack_11937_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 165_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_K9_13851_delayed_9_13910_inst_ack_0, ack => e_block_daemon_CP_11105_elements(165)); -- 
    -- CP-element group 166:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	164 
    -- CP-element group 166: successors 
    -- CP-element group 166: 	167 
    -- CP-element group 166: marked-successors 
    -- CP-element group 166: 	164 
    -- CP-element group 166:  members (7) 
      -- CP-element group 166: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13912_update_completed_
      -- CP-element group 166: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13912_Update/$exit
      -- CP-element group 166: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13912_Update/ack
      -- CP-element group 166: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_K9_13851_delayed_9_13914_sample_start_
      -- CP-element group 166: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_K9_13851_delayed_9_13914_sample_completed_
      -- CP-element group 166: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_K9_13851_delayed_9_13914_update_start_
      -- CP-element group 166: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_K9_13851_delayed_9_13914_update_completed_
      -- 
    ack_11942_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 166_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_K9_13851_delayed_9_13910_inst_ack_1, ack => e_block_daemon_CP_11105_elements(166)); -- 
    -- CP-element group 167:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	161 
    -- CP-element group 167: 	166 
    -- CP-element group 167: marked-predecessors 
    -- CP-element group 167: 	169 
    -- CP-element group 167: successors 
    -- CP-element group 167: 	169 
    -- CP-element group 167:  members (3) 
      -- CP-element group 167: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13917_sample_start_
      -- CP-element group 167: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13917_Sample/$entry
      -- CP-element group 167: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13917_Sample/crr
      -- 
    crr_11958_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_11958_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_block_daemon_CP_11105_elements(167), ack => call_stmt_13917_call_req_0); -- 
    e_block_daemon_cp_element_group_167: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 2,1 => 2,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 35) := "e_block_daemon_cp_element_group_167"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= e_block_daemon_CP_11105_elements(161) & e_block_daemon_CP_11105_elements(166) & e_block_daemon_CP_11105_elements(169);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => e_block_daemon_CP_11105_elements(167), clk => clk, reset => reset); --
    end block;
    -- CP-element group 168:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	58 
    -- CP-element group 168: marked-predecessors 
    -- CP-element group 168: 	170 
    -- CP-element group 168: 	178 
    -- CP-element group 168: successors 
    -- CP-element group 168: 	170 
    -- CP-element group 168:  members (3) 
      -- CP-element group 168: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13917_update_start_
      -- CP-element group 168: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13917_Update/$entry
      -- CP-element group 168: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13917_Update/ccr
      -- 
    ccr_11963_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_11963_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_block_daemon_CP_11105_elements(168), ack => call_stmt_13917_call_req_1); -- 
    e_block_daemon_cp_element_group_168: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 2,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "e_block_daemon_cp_element_group_168"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= e_block_daemon_CP_11105_elements(58) & e_block_daemon_CP_11105_elements(170) & e_block_daemon_CP_11105_elements(178);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => e_block_daemon_CP_11105_elements(168), clk => clk, reset => reset); --
    end block;
    -- CP-element group 169:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	167 
    -- CP-element group 169: successors 
    -- CP-element group 169: marked-successors 
    -- CP-element group 169: 	159 
    -- CP-element group 169: 	164 
    -- CP-element group 169: 	167 
    -- CP-element group 169:  members (3) 
      -- CP-element group 169: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13917_sample_completed_
      -- CP-element group 169: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13917_Sample/$exit
      -- CP-element group 169: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13917_Sample/cra
      -- 
    cra_11959_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 169_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_13917_call_ack_0, ack => e_block_daemon_CP_11105_elements(169)); -- 
    -- CP-element group 170:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	168 
    -- CP-element group 170: successors 
    -- CP-element group 170: 	176 
    -- CP-element group 170: marked-successors 
    -- CP-element group 170: 	168 
    -- CP-element group 170:  members (7) 
      -- CP-element group 170: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13917_update_completed_
      -- CP-element group 170: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13917_Update/$exit
      -- CP-element group 170: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13917_Update/cca
      -- CP-element group 170: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_round_S9_13921_sample_start_
      -- CP-element group 170: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_round_S9_13921_sample_completed_
      -- CP-element group 170: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_round_S9_13921_update_start_
      -- CP-element group 170: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_round_S9_13921_update_completed_
      -- 
    cca_11964_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 170_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_13917_call_ack_1, ack => e_block_daemon_CP_11105_elements(170)); -- 
    -- CP-element group 171:  join  transition  bypass  pipeline-parent 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	58 
    -- CP-element group 171: marked-predecessors 
    -- CP-element group 171: 	174 
    -- CP-element group 171: successors 
    -- CP-element group 171: 	172 
    -- CP-element group 171:  members (2) 
      -- CP-element group 171: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_K10_13919_update_start_
      -- CP-element group 171: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_K10_13919_update_completed_
      -- 
    e_block_daemon_cp_element_group_171: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 2,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "e_block_daemon_cp_element_group_171"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= e_block_daemon_CP_11105_elements(58) & e_block_daemon_CP_11105_elements(174);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => e_block_daemon_CP_11105_elements(171), clk => clk, reset => reset); --
    end block;
    -- CP-element group 172:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	171 
    -- CP-element group 172: marked-predecessors 
    -- CP-element group 172: 	174 
    -- CP-element group 172: successors 
    -- CP-element group 172: 	174 
    -- CP-element group 172:  members (3) 
      -- CP-element group 172: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13920_sample_start_
      -- CP-element group 172: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13920_Sample/$entry
      -- CP-element group 172: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13920_Sample/req
      -- 
    req_11976_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_11976_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_block_daemon_CP_11105_elements(172), ack => W_K10_13856_delayed_10_13918_inst_req_0); -- 
    e_block_daemon_cp_element_group_172: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 2,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "e_block_daemon_cp_element_group_172"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= e_block_daemon_CP_11105_elements(171) & e_block_daemon_CP_11105_elements(174);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => e_block_daemon_CP_11105_elements(172), clk => clk, reset => reset); --
    end block;
    -- CP-element group 173:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	58 
    -- CP-element group 173: marked-predecessors 
    -- CP-element group 173: 	175 
    -- CP-element group 173: 	178 
    -- CP-element group 173: successors 
    -- CP-element group 173: 	175 
    -- CP-element group 173:  members (3) 
      -- CP-element group 173: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13920_update_start_
      -- CP-element group 173: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13920_Update/$entry
      -- CP-element group 173: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13920_Update/req
      -- 
    req_11981_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_11981_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_block_daemon_CP_11105_elements(173), ack => W_K10_13856_delayed_10_13918_inst_req_1); -- 
    e_block_daemon_cp_element_group_173: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 2,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "e_block_daemon_cp_element_group_173"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= e_block_daemon_CP_11105_elements(58) & e_block_daemon_CP_11105_elements(175) & e_block_daemon_CP_11105_elements(178);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => e_block_daemon_CP_11105_elements(173), clk => clk, reset => reset); --
    end block;
    -- CP-element group 174:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	172 
    -- CP-element group 174: successors 
    -- CP-element group 174: marked-successors 
    -- CP-element group 174: 	171 
    -- CP-element group 174: 	172 
    -- CP-element group 174:  members (3) 
      -- CP-element group 174: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13920_sample_completed_
      -- CP-element group 174: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13920_Sample/$exit
      -- CP-element group 174: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13920_Sample/ack
      -- 
    ack_11977_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 174_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_K10_13856_delayed_10_13918_inst_ack_0, ack => e_block_daemon_CP_11105_elements(174)); -- 
    -- CP-element group 175:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	173 
    -- CP-element group 175: successors 
    -- CP-element group 175: 	176 
    -- CP-element group 175: marked-successors 
    -- CP-element group 175: 	173 
    -- CP-element group 175:  members (7) 
      -- CP-element group 175: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13920_update_completed_
      -- CP-element group 175: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13920_Update/$exit
      -- CP-element group 175: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/assign_stmt_13920_Update/ack
      -- CP-element group 175: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_K10_13856_delayed_10_13922_sample_start_
      -- CP-element group 175: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_K10_13856_delayed_10_13922_sample_completed_
      -- CP-element group 175: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_K10_13856_delayed_10_13922_update_start_
      -- CP-element group 175: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_K10_13856_delayed_10_13922_update_completed_
      -- 
    ack_11982_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 175_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_K10_13856_delayed_10_13918_inst_ack_1, ack => e_block_daemon_CP_11105_elements(175)); -- 
    -- CP-element group 176:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: 	170 
    -- CP-element group 176: 	175 
    -- CP-element group 176: marked-predecessors 
    -- CP-element group 176: 	178 
    -- CP-element group 176: successors 
    -- CP-element group 176: 	178 
    -- CP-element group 176:  members (3) 
      -- CP-element group 176: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13925_sample_start_
      -- CP-element group 176: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13925_Sample/$entry
      -- CP-element group 176: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13925_Sample/crr
      -- 
    crr_11998_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_11998_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_block_daemon_CP_11105_elements(176), ack => call_stmt_13925_call_req_0); -- 
    e_block_daemon_cp_element_group_176: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 2,1 => 2,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 35) := "e_block_daemon_cp_element_group_176"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= e_block_daemon_CP_11105_elements(170) & e_block_daemon_CP_11105_elements(175) & e_block_daemon_CP_11105_elements(178);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => e_block_daemon_CP_11105_elements(176), clk => clk, reset => reset); --
    end block;
    -- CP-element group 177:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	58 
    -- CP-element group 177: marked-predecessors 
    -- CP-element group 177: 	179 
    -- CP-element group 177: 	182 
    -- CP-element group 177: successors 
    -- CP-element group 177: 	179 
    -- CP-element group 177:  members (3) 
      -- CP-element group 177: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13925_update_start_
      -- CP-element group 177: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13925_Update/$entry
      -- CP-element group 177: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13925_Update/ccr
      -- 
    ccr_12003_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_12003_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_block_daemon_CP_11105_elements(177), ack => call_stmt_13925_call_req_1); -- 
    e_block_daemon_cp_element_group_177: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 2,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "e_block_daemon_cp_element_group_177"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= e_block_daemon_CP_11105_elements(58) & e_block_daemon_CP_11105_elements(179) & e_block_daemon_CP_11105_elements(182);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => e_block_daemon_CP_11105_elements(177), clk => clk, reset => reset); --
    end block;
    -- CP-element group 178:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	176 
    -- CP-element group 178: successors 
    -- CP-element group 178: marked-successors 
    -- CP-element group 178: 	168 
    -- CP-element group 178: 	173 
    -- CP-element group 178: 	176 
    -- CP-element group 178:  members (3) 
      -- CP-element group 178: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13925_sample_completed_
      -- CP-element group 178: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13925_Sample/$exit
      -- CP-element group 178: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13925_Sample/cra
      -- 
    cra_11999_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 178_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_13925_call_ack_0, ack => e_block_daemon_CP_11105_elements(178)); -- 
    -- CP-element group 179:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	177 
    -- CP-element group 179: successors 
    -- CP-element group 179: 	180 
    -- CP-element group 179: marked-successors 
    -- CP-element group 179: 	177 
    -- CP-element group 179:  members (7) 
      -- CP-element group 179: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13925_update_completed_
      -- CP-element group 179: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13925_Update/$exit
      -- CP-element group 179: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/call_stmt_13925_Update/cca
      -- CP-element group 179: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_round_S10_13927_sample_start_
      -- CP-element group 179: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_round_S10_13927_sample_completed_
      -- CP-element group 179: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_round_S10_13927_update_start_
      -- CP-element group 179: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_round_S10_13927_update_completed_
      -- 
    cca_12004_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 179_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_13925_call_ack_1, ack => e_block_daemon_CP_11105_elements(179)); -- 
    -- CP-element group 180:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	179 
    -- CP-element group 180: marked-predecessors 
    -- CP-element group 180: 	182 
    -- CP-element group 180: successors 
    -- CP-element group 180: 	182 
    -- CP-element group 180:  members (3) 
      -- CP-element group 180: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/WPIPE_e_out_buf_13926_sample_start_
      -- CP-element group 180: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/WPIPE_e_out_buf_13926_Sample/$entry
      -- CP-element group 180: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/WPIPE_e_out_buf_13926_Sample/req
      -- 
    req_12016_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_12016_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_block_daemon_CP_11105_elements(180), ack => WPIPE_e_out_buf_13926_inst_req_0); -- 
    e_block_daemon_cp_element_group_180: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 2,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "e_block_daemon_cp_element_group_180"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= e_block_daemon_CP_11105_elements(179) & e_block_daemon_CP_11105_elements(182);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => e_block_daemon_CP_11105_elements(180), clk => clk, reset => reset); --
    end block;
    -- CP-element group 181:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	182 
    -- CP-element group 181: marked-predecessors 
    -- CP-element group 181: 	183 
    -- CP-element group 181: successors 
    -- CP-element group 181: 	183 
    -- CP-element group 181:  members (3) 
      -- CP-element group 181: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/WPIPE_e_out_buf_13926_update_start_
      -- CP-element group 181: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/WPIPE_e_out_buf_13926_Update/$entry
      -- CP-element group 181: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/WPIPE_e_out_buf_13926_Update/req
      -- 
    req_12021_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_12021_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_block_daemon_CP_11105_elements(181), ack => WPIPE_e_out_buf_13926_inst_req_1); -- 
    e_block_daemon_cp_element_group_181: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 2,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "e_block_daemon_cp_element_group_181"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= e_block_daemon_CP_11105_elements(182) & e_block_daemon_CP_11105_elements(183);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => e_block_daemon_CP_11105_elements(181), clk => clk, reset => reset); --
    end block;
    -- CP-element group 182:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	180 
    -- CP-element group 182: successors 
    -- CP-element group 182: 	181 
    -- CP-element group 182: marked-successors 
    -- CP-element group 182: 	177 
    -- CP-element group 182: 	180 
    -- CP-element group 182:  members (3) 
      -- CP-element group 182: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/WPIPE_e_out_buf_13926_sample_completed_
      -- CP-element group 182: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/WPIPE_e_out_buf_13926_Sample/$exit
      -- CP-element group 182: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/WPIPE_e_out_buf_13926_Sample/ack
      -- 
    ack_12017_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 182_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_e_out_buf_13926_inst_ack_0, ack => e_block_daemon_CP_11105_elements(182)); -- 
    -- CP-element group 183:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: 	181 
    -- CP-element group 183: successors 
    -- CP-element group 183: 	249 
    -- CP-element group 183: marked-successors 
    -- CP-element group 183: 	181 
    -- CP-element group 183:  members (3) 
      -- CP-element group 183: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/WPIPE_e_out_buf_13926_update_completed_
      -- CP-element group 183: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/WPIPE_e_out_buf_13926_Update/$exit
      -- CP-element group 183: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/WPIPE_e_out_buf_13926_Update/ack
      -- 
    ack_12022_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 183_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_e_out_buf_13926_inst_ack_1, ack => e_block_daemon_CP_11105_elements(183)); -- 
    -- CP-element group 184:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	63 
    -- CP-element group 184: marked-predecessors 
    -- CP-element group 184: 	186 
    -- CP-element group 184: successors 
    -- CP-element group 184: 	186 
    -- CP-element group 184:  members (3) 
      -- CP-element group 184: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/ADD_u15_u15_13932_sample_start_
      -- CP-element group 184: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/ADD_u15_u15_13932_Sample/$entry
      -- CP-element group 184: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/ADD_u15_u15_13932_Sample/rr
      -- 
    rr_12034_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_12034_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_block_daemon_CP_11105_elements(184), ack => ADD_u15_u15_13932_inst_req_0); -- 
    e_block_daemon_cp_element_group_184: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 2,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "e_block_daemon_cp_element_group_184"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= e_block_daemon_CP_11105_elements(63) & e_block_daemon_CP_11105_elements(186);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => e_block_daemon_CP_11105_elements(184), clk => clk, reset => reset); --
    end block;
    -- CP-element group 185:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	62 
    -- CP-element group 185: marked-predecessors 
    -- CP-element group 185: 	187 
    -- CP-element group 185: successors 
    -- CP-element group 185: 	187 
    -- CP-element group 185:  members (3) 
      -- CP-element group 185: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/ADD_u15_u15_13932_update_start_
      -- CP-element group 185: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/ADD_u15_u15_13932_Update/$entry
      -- CP-element group 185: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/ADD_u15_u15_13932_Update/cr
      -- 
    cr_12039_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_12039_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_block_daemon_CP_11105_elements(185), ack => ADD_u15_u15_13932_inst_req_1); -- 
    e_block_daemon_cp_element_group_185: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 2,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "e_block_daemon_cp_element_group_185"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= e_block_daemon_CP_11105_elements(62) & e_block_daemon_CP_11105_elements(187);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => e_block_daemon_CP_11105_elements(185), clk => clk, reset => reset); --
    end block;
    -- CP-element group 186:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	184 
    -- CP-element group 186: successors 
    -- CP-element group 186: marked-successors 
    -- CP-element group 186: 	184 
    -- CP-element group 186: 	61 
    -- CP-element group 186:  members (3) 
      -- CP-element group 186: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/ADD_u15_u15_13932_sample_completed_
      -- CP-element group 186: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/ADD_u15_u15_13932_Sample/$exit
      -- CP-element group 186: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/ADD_u15_u15_13932_Sample/ra
      -- 
    ra_12035_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 186_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u15_u15_13932_inst_ack_0, ack => e_block_daemon_CP_11105_elements(186)); -- 
    -- CP-element group 187:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: 	185 
    -- CP-element group 187: successors 
    -- CP-element group 187: 	188 
    -- CP-element group 187: marked-successors 
    -- CP-element group 187: 	185 
    -- CP-element group 187: 	60 
    -- CP-element group 187:  members (7) 
      -- CP-element group 187: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/ADD_u15_u15_13932_update_completed_
      -- CP-element group 187: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/ADD_u15_u15_13932_Update/$exit
      -- CP-element group 187: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/ADD_u15_u15_13932_Update/ca
      -- CP-element group 187: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_n_count_var_13935_sample_start_
      -- CP-element group 187: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_n_count_var_13935_sample_completed_
      -- CP-element group 187: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_n_count_var_13935_update_start_
      -- CP-element group 187: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/R_n_count_var_13935_update_completed_
      -- 
    ca_12040_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 187_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u15_u15_13932_inst_ack_1, ack => e_block_daemon_CP_11105_elements(187)); -- 
    -- CP-element group 188:  join  transition  bypass  pipeline-parent 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: 	187 
    -- CP-element group 188: 	58 
    -- CP-element group 188: successors 
    -- CP-element group 188: 	59 
    -- CP-element group 188:  members (12) 
      -- CP-element group 188: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/ULT_u15_u1_13937_sample_start_
      -- CP-element group 188: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/ULT_u15_u1_13937_sample_completed_
      -- CP-element group 188: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/ULT_u15_u1_13937_update_start_
      -- CP-element group 188: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/ULT_u15_u1_13937_update_completed_
      -- CP-element group 188: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/ULT_u15_u1_13937_Sample/$entry
      -- CP-element group 188: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/ULT_u15_u1_13937_Sample/$exit
      -- CP-element group 188: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/ULT_u15_u1_13937_Sample/rr
      -- CP-element group 188: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/ULT_u15_u1_13937_Sample/ra
      -- CP-element group 188: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/ULT_u15_u1_13937_Update/$entry
      -- CP-element group 188: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/ULT_u15_u1_13937_Update/$exit
      -- CP-element group 188: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/ULT_u15_u1_13937_Update/cr
      -- CP-element group 188: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/ULT_u15_u1_13937_Update/ca
      -- 
    e_block_daemon_cp_element_group_188: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 2,1 => 2);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "e_block_daemon_cp_element_group_188"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= e_block_daemon_CP_11105_elements(187) & e_block_daemon_CP_11105_elements(58);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => e_block_daemon_CP_11105_elements(188), clk => clk, reset => reset); --
    end block;
    -- CP-element group 189:  transition  bypass  pipeline-parent 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: 	54 
    -- CP-element group 189: successors 
    -- CP-element group 189: 	190 
    -- CP-element group 189:  members (1) 
      -- CP-element group 189: 	 branch_block_stmt_13736/do_while_stmt_13828/loop_exit/$entry
      -- 
    e_block_daemon_CP_11105_elements(189) <= e_block_daemon_CP_11105_elements(54);
    -- CP-element group 190:  transition  input  bypass  pipeline-parent 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: 	189 
    -- CP-element group 190: successors 
    -- CP-element group 190:  members (2) 
      -- CP-element group 190: 	 branch_block_stmt_13736/do_while_stmt_13828/loop_exit/$exit
      -- CP-element group 190: 	 branch_block_stmt_13736/do_while_stmt_13828/loop_exit/ack
      -- 
    ack_12066_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 190_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_13828_branch_ack_0, ack => e_block_daemon_CP_11105_elements(190)); -- 
    -- CP-element group 191:  transition  bypass  pipeline-parent 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: 	54 
    -- CP-element group 191: successors 
    -- CP-element group 191: 	192 
    -- CP-element group 191:  members (1) 
      -- CP-element group 191: 	 branch_block_stmt_13736/do_while_stmt_13828/loop_taken/$entry
      -- 
    e_block_daemon_CP_11105_elements(191) <= e_block_daemon_CP_11105_elements(54);
    -- CP-element group 192:  transition  input  bypass  pipeline-parent 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: 	191 
    -- CP-element group 192: successors 
    -- CP-element group 192:  members (2) 
      -- CP-element group 192: 	 branch_block_stmt_13736/do_while_stmt_13828/loop_taken/$exit
      -- CP-element group 192: 	 branch_block_stmt_13736/do_while_stmt_13828/loop_taken/ack
      -- 
    ack_12070_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 192_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_13828_branch_ack_1, ack => e_block_daemon_CP_11105_elements(192)); -- 
    -- CP-element group 193:  transition  bypass  pipeline-parent 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: 	52 
    -- CP-element group 193: successors 
    -- CP-element group 193: 	10 
    -- CP-element group 193:  members (1) 
      -- CP-element group 193: 	 branch_block_stmt_13736/do_while_stmt_13828/$exit
      -- 
    e_block_daemon_CP_11105_elements(193) <= e_block_daemon_CP_11105_elements(52);
    -- CP-element group 194:  transition  output  bypass 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: 	10 
    -- CP-element group 194: successors 
    -- CP-element group 194: 	195 
    -- CP-element group 194:  members (4) 
      -- CP-element group 194: 	 branch_block_stmt_13736/assign_stmt_13940/$entry
      -- CP-element group 194: 	 branch_block_stmt_13736/assign_stmt_13940/WPIPE_e_block_done_13938_sample_start_
      -- CP-element group 194: 	 branch_block_stmt_13736/assign_stmt_13940/WPIPE_e_block_done_13938_Sample/$entry
      -- CP-element group 194: 	 branch_block_stmt_13736/assign_stmt_13940/WPIPE_e_block_done_13938_Sample/req
      -- 
    req_12082_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_12082_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_block_daemon_CP_11105_elements(194), ack => WPIPE_e_block_done_13938_inst_req_0); -- 
    e_block_daemon_CP_11105_elements(194) <= e_block_daemon_CP_11105_elements(10);
    -- CP-element group 195:  transition  input  output  bypass 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: 	194 
    -- CP-element group 195: successors 
    -- CP-element group 195: 	196 
    -- CP-element group 195:  members (6) 
      -- CP-element group 195: 	 branch_block_stmt_13736/assign_stmt_13940/WPIPE_e_block_done_13938_sample_completed_
      -- CP-element group 195: 	 branch_block_stmt_13736/assign_stmt_13940/WPIPE_e_block_done_13938_update_start_
      -- CP-element group 195: 	 branch_block_stmt_13736/assign_stmt_13940/WPIPE_e_block_done_13938_Sample/$exit
      -- CP-element group 195: 	 branch_block_stmt_13736/assign_stmt_13940/WPIPE_e_block_done_13938_Sample/ack
      -- CP-element group 195: 	 branch_block_stmt_13736/assign_stmt_13940/WPIPE_e_block_done_13938_Update/$entry
      -- CP-element group 195: 	 branch_block_stmt_13736/assign_stmt_13940/WPIPE_e_block_done_13938_Update/req
      -- 
    ack_12083_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 195_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_e_block_done_13938_inst_ack_0, ack => e_block_daemon_CP_11105_elements(195)); -- 
    req_12087_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_12087_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_block_daemon_CP_11105_elements(195), ack => WPIPE_e_block_done_13938_inst_req_1); -- 
    -- CP-element group 196:  transition  input  bypass 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: 	195 
    -- CP-element group 196: successors 
    -- CP-element group 196: 	11 
    -- CP-element group 196:  members (4) 
      -- CP-element group 196: 	 branch_block_stmt_13736/assign_stmt_13940/$exit
      -- CP-element group 196: 	 branch_block_stmt_13736/assign_stmt_13940/WPIPE_e_block_done_13938_update_completed_
      -- CP-element group 196: 	 branch_block_stmt_13736/assign_stmt_13940/WPIPE_e_block_done_13938_Update/$exit
      -- CP-element group 196: 	 branch_block_stmt_13736/assign_stmt_13940/WPIPE_e_block_done_13938_Update/ack
      -- 
    ack_12088_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 196_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_e_block_done_13938_inst_ack_1, ack => e_block_daemon_CP_11105_elements(196)); -- 
    -- CP-element group 197:  transition  output  bypass 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: 	11 
    -- CP-element group 197: successors 
    -- CP-element group 197: 	198 
    -- CP-element group 197:  members (4) 
      -- CP-element group 197: 	 branch_block_stmt_13736/assign_stmt_13943/$entry
      -- CP-element group 197: 	 branch_block_stmt_13736/assign_stmt_13943/RPIPE_e_cmd_pipe_13942_sample_start_
      -- CP-element group 197: 	 branch_block_stmt_13736/assign_stmt_13943/RPIPE_e_cmd_pipe_13942_Sample/$entry
      -- CP-element group 197: 	 branch_block_stmt_13736/assign_stmt_13943/RPIPE_e_cmd_pipe_13942_Sample/rr
      -- 
    rr_12099_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_12099_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_block_daemon_CP_11105_elements(197), ack => RPIPE_e_cmd_pipe_13942_inst_req_0); -- 
    e_block_daemon_CP_11105_elements(197) <= e_block_daemon_CP_11105_elements(11);
    -- CP-element group 198:  transition  input  output  bypass 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: 	197 
    -- CP-element group 198: successors 
    -- CP-element group 198: 	199 
    -- CP-element group 198:  members (6) 
      -- CP-element group 198: 	 branch_block_stmt_13736/assign_stmt_13943/RPIPE_e_cmd_pipe_13942_sample_completed_
      -- CP-element group 198: 	 branch_block_stmt_13736/assign_stmt_13943/RPIPE_e_cmd_pipe_13942_update_start_
      -- CP-element group 198: 	 branch_block_stmt_13736/assign_stmt_13943/RPIPE_e_cmd_pipe_13942_Sample/$exit
      -- CP-element group 198: 	 branch_block_stmt_13736/assign_stmt_13943/RPIPE_e_cmd_pipe_13942_Sample/ra
      -- CP-element group 198: 	 branch_block_stmt_13736/assign_stmt_13943/RPIPE_e_cmd_pipe_13942_Update/$entry
      -- CP-element group 198: 	 branch_block_stmt_13736/assign_stmt_13943/RPIPE_e_cmd_pipe_13942_Update/cr
      -- 
    ra_12100_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 198_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_e_cmd_pipe_13942_inst_ack_0, ack => e_block_daemon_CP_11105_elements(198)); -- 
    cr_12104_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_12104_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_block_daemon_CP_11105_elements(198), ack => RPIPE_e_cmd_pipe_13942_inst_req_1); -- 
    -- CP-element group 199:  transition  input  bypass 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: 	198 
    -- CP-element group 199: successors 
    -- CP-element group 199: 	12 
    -- CP-element group 199:  members (4) 
      -- CP-element group 199: 	 branch_block_stmt_13736/assign_stmt_13943/$exit
      -- CP-element group 199: 	 branch_block_stmt_13736/assign_stmt_13943/RPIPE_e_cmd_pipe_13942_update_completed_
      -- CP-element group 199: 	 branch_block_stmt_13736/assign_stmt_13943/RPIPE_e_cmd_pipe_13942_Update/$exit
      -- CP-element group 199: 	 branch_block_stmt_13736/assign_stmt_13943/RPIPE_e_cmd_pipe_13942_Update/ca
      -- 
    ca_12105_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 199_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_e_cmd_pipe_13942_inst_ack_1, ack => e_block_daemon_CP_11105_elements(199)); -- 
    -- CP-element group 200:  join  fork  transition  bypass 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: 	12 
    -- CP-element group 200: successors 
    -- CP-element group 200: 	13 
    -- CP-element group 200:  members (50) 
      -- CP-element group 200: 	 branch_block_stmt_13736/assign_stmt_13947_to_assign_stmt_13955/slice_13954_Update/cr
      -- CP-element group 200: 	 branch_block_stmt_13736/assign_stmt_13947_to_assign_stmt_13955/slice_13954_Update/$entry
      -- CP-element group 200: 	 branch_block_stmt_13736/assign_stmt_13947_to_assign_stmt_13955/slice_13954_Update/$exit
      -- CP-element group 200: 	 branch_block_stmt_13736/assign_stmt_13947_to_assign_stmt_13955/slice_13954_Update/ca
      -- CP-element group 200: 	 branch_block_stmt_13736/assign_stmt_13947_to_assign_stmt_13955/$entry
      -- CP-element group 200: 	 branch_block_stmt_13736/assign_stmt_13947_to_assign_stmt_13955/$exit
      -- CP-element group 200: 	 branch_block_stmt_13736/assign_stmt_13947_to_assign_stmt_13955/slice_13946_sample_start_
      -- CP-element group 200: 	 branch_block_stmt_13736/assign_stmt_13947_to_assign_stmt_13955/slice_13946_sample_completed_
      -- CP-element group 200: 	 branch_block_stmt_13736/assign_stmt_13947_to_assign_stmt_13955/slice_13946_update_start_
      -- CP-element group 200: 	 branch_block_stmt_13736/assign_stmt_13947_to_assign_stmt_13955/slice_13946_update_completed_
      -- CP-element group 200: 	 branch_block_stmt_13736/assign_stmt_13947_to_assign_stmt_13955/R_e_new_cmd_13945_sample_start_
      -- CP-element group 200: 	 branch_block_stmt_13736/assign_stmt_13947_to_assign_stmt_13955/R_e_new_cmd_13945_sample_completed_
      -- CP-element group 200: 	 branch_block_stmt_13736/assign_stmt_13947_to_assign_stmt_13955/R_e_new_cmd_13945_update_start_
      -- CP-element group 200: 	 branch_block_stmt_13736/assign_stmt_13947_to_assign_stmt_13955/R_e_new_cmd_13945_update_completed_
      -- CP-element group 200: 	 branch_block_stmt_13736/assign_stmt_13947_to_assign_stmt_13955/slice_13946_Sample/$entry
      -- CP-element group 200: 	 branch_block_stmt_13736/assign_stmt_13947_to_assign_stmt_13955/slice_13946_Sample/$exit
      -- CP-element group 200: 	 branch_block_stmt_13736/assign_stmt_13947_to_assign_stmt_13955/slice_13946_Sample/rr
      -- CP-element group 200: 	 branch_block_stmt_13736/assign_stmt_13947_to_assign_stmt_13955/slice_13946_Sample/ra
      -- CP-element group 200: 	 branch_block_stmt_13736/assign_stmt_13947_to_assign_stmt_13955/slice_13946_Update/$entry
      -- CP-element group 200: 	 branch_block_stmt_13736/assign_stmt_13947_to_assign_stmt_13955/slice_13946_Update/$exit
      -- CP-element group 200: 	 branch_block_stmt_13736/assign_stmt_13947_to_assign_stmt_13955/slice_13946_Update/cr
      -- CP-element group 200: 	 branch_block_stmt_13736/assign_stmt_13947_to_assign_stmt_13955/slice_13946_Update/ca
      -- CP-element group 200: 	 branch_block_stmt_13736/assign_stmt_13947_to_assign_stmt_13955/slice_13950_sample_start_
      -- CP-element group 200: 	 branch_block_stmt_13736/assign_stmt_13947_to_assign_stmt_13955/slice_13950_sample_completed_
      -- CP-element group 200: 	 branch_block_stmt_13736/assign_stmt_13947_to_assign_stmt_13955/slice_13950_update_start_
      -- CP-element group 200: 	 branch_block_stmt_13736/assign_stmt_13947_to_assign_stmt_13955/slice_13950_update_completed_
      -- CP-element group 200: 	 branch_block_stmt_13736/assign_stmt_13947_to_assign_stmt_13955/R_e_new_cmd_13949_sample_start_
      -- CP-element group 200: 	 branch_block_stmt_13736/assign_stmt_13947_to_assign_stmt_13955/R_e_new_cmd_13949_sample_completed_
      -- CP-element group 200: 	 branch_block_stmt_13736/assign_stmt_13947_to_assign_stmt_13955/R_e_new_cmd_13949_update_start_
      -- CP-element group 200: 	 branch_block_stmt_13736/assign_stmt_13947_to_assign_stmt_13955/R_e_new_cmd_13949_update_completed_
      -- CP-element group 200: 	 branch_block_stmt_13736/assign_stmt_13947_to_assign_stmt_13955/slice_13950_Sample/$entry
      -- CP-element group 200: 	 branch_block_stmt_13736/assign_stmt_13947_to_assign_stmt_13955/slice_13950_Sample/$exit
      -- CP-element group 200: 	 branch_block_stmt_13736/assign_stmt_13947_to_assign_stmt_13955/slice_13950_Sample/rr
      -- CP-element group 200: 	 branch_block_stmt_13736/assign_stmt_13947_to_assign_stmt_13955/slice_13950_Sample/ra
      -- CP-element group 200: 	 branch_block_stmt_13736/assign_stmt_13947_to_assign_stmt_13955/slice_13950_Update/$entry
      -- CP-element group 200: 	 branch_block_stmt_13736/assign_stmt_13947_to_assign_stmt_13955/slice_13950_Update/$exit
      -- CP-element group 200: 	 branch_block_stmt_13736/assign_stmt_13947_to_assign_stmt_13955/slice_13950_Update/cr
      -- CP-element group 200: 	 branch_block_stmt_13736/assign_stmt_13947_to_assign_stmt_13955/slice_13950_Update/ca
      -- CP-element group 200: 	 branch_block_stmt_13736/assign_stmt_13947_to_assign_stmt_13955/slice_13954_sample_start_
      -- CP-element group 200: 	 branch_block_stmt_13736/assign_stmt_13947_to_assign_stmt_13955/slice_13954_sample_completed_
      -- CP-element group 200: 	 branch_block_stmt_13736/assign_stmt_13947_to_assign_stmt_13955/slice_13954_update_start_
      -- CP-element group 200: 	 branch_block_stmt_13736/assign_stmt_13947_to_assign_stmt_13955/slice_13954_update_completed_
      -- CP-element group 200: 	 branch_block_stmt_13736/assign_stmt_13947_to_assign_stmt_13955/R_e_new_cmd_13953_sample_start_
      -- CP-element group 200: 	 branch_block_stmt_13736/assign_stmt_13947_to_assign_stmt_13955/R_e_new_cmd_13953_sample_completed_
      -- CP-element group 200: 	 branch_block_stmt_13736/assign_stmt_13947_to_assign_stmt_13955/R_e_new_cmd_13953_update_start_
      -- CP-element group 200: 	 branch_block_stmt_13736/assign_stmt_13947_to_assign_stmt_13955/R_e_new_cmd_13953_update_completed_
      -- CP-element group 200: 	 branch_block_stmt_13736/assign_stmt_13947_to_assign_stmt_13955/slice_13954_Sample/$entry
      -- CP-element group 200: 	 branch_block_stmt_13736/assign_stmt_13947_to_assign_stmt_13955/slice_13954_Sample/$exit
      -- CP-element group 200: 	 branch_block_stmt_13736/assign_stmt_13947_to_assign_stmt_13955/slice_13954_Sample/rr
      -- CP-element group 200: 	 branch_block_stmt_13736/assign_stmt_13947_to_assign_stmt_13955/slice_13954_Sample/ra
      -- 
    e_block_daemon_CP_11105_elements(200) <= e_block_daemon_CP_11105_elements(12);
    -- CP-element group 201:  transition  bypass 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: 	13 
    -- CP-element group 201: successors 
    -- CP-element group 201:  members (1) 
      -- CP-element group 201: 	 branch_block_stmt_13736/if_stmt_13956_dead_link/$entry
      -- 
    e_block_daemon_CP_11105_elements(201) <= e_block_daemon_CP_11105_elements(13);
    -- CP-element group 202:  transition  output  bypass 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: 	13 
    -- CP-element group 202: successors 
    -- CP-element group 202: 	203 
    -- CP-element group 202:  members (17) 
      -- CP-element group 202: 	 branch_block_stmt_13736/if_stmt_13956_eval_test/EQ_u1_u1_13959/$entry
      -- CP-element group 202: 	 branch_block_stmt_13736/if_stmt_13956_eval_test/$exit
      -- CP-element group 202: 	 branch_block_stmt_13736/if_stmt_13956_eval_test/EQ_u1_u1_13959/EQ_u1_u1_13959_inputs/$exit
      -- CP-element group 202: 	 branch_block_stmt_13736/if_stmt_13956_eval_test/EQ_u1_u1_13959/EQ_u1_u1_13959_inputs/$entry
      -- CP-element group 202: 	 branch_block_stmt_13736/if_stmt_13956_eval_test/$entry
      -- CP-element group 202: 	 branch_block_stmt_13736/if_stmt_13956_eval_test/EQ_u1_u1_13959/SplitProtocol/$entry
      -- CP-element group 202: 	 branch_block_stmt_13736/if_stmt_13956_eval_test/branch_req
      -- CP-element group 202: 	 branch_block_stmt_13736/if_stmt_13956_eval_test/EQ_u1_u1_13959/SplitProtocol/Update/ca
      -- CP-element group 202: 	 branch_block_stmt_13736/if_stmt_13956_eval_test/EQ_u1_u1_13959/SplitProtocol/Update/cr
      -- CP-element group 202: 	 branch_block_stmt_13736/if_stmt_13956_eval_test/EQ_u1_u1_13959/SplitProtocol/Update/$exit
      -- CP-element group 202: 	 branch_block_stmt_13736/if_stmt_13956_eval_test/EQ_u1_u1_13959/SplitProtocol/Update/$entry
      -- CP-element group 202: 	 branch_block_stmt_13736/if_stmt_13956_eval_test/EQ_u1_u1_13959/SplitProtocol/Sample/ra
      -- CP-element group 202: 	 branch_block_stmt_13736/if_stmt_13956_eval_test/EQ_u1_u1_13959/SplitProtocol/Sample/rr
      -- CP-element group 202: 	 branch_block_stmt_13736/if_stmt_13956_eval_test/EQ_u1_u1_13959/SplitProtocol/Sample/$exit
      -- CP-element group 202: 	 branch_block_stmt_13736/if_stmt_13956_eval_test/EQ_u1_u1_13959/SplitProtocol/Sample/$entry
      -- CP-element group 202: 	 branch_block_stmt_13736/if_stmt_13956_eval_test/EQ_u1_u1_13959/SplitProtocol/$exit
      -- CP-element group 202: 	 branch_block_stmt_13736/if_stmt_13956_eval_test/EQ_u1_u1_13959/$exit
      -- 
    branch_req_12189_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_12189_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_block_daemon_CP_11105_elements(202), ack => if_stmt_13956_branch_req_0); -- 
    e_block_daemon_CP_11105_elements(202) <= e_block_daemon_CP_11105_elements(13);
    -- CP-element group 203:  branch  place  bypass 
    -- CP-element group 203: predecessors 
    -- CP-element group 203: 	202 
    -- CP-element group 203: successors 
    -- CP-element group 203: 	204 
    -- CP-element group 203: 	206 
    -- CP-element group 203:  members (1) 
      -- CP-element group 203: 	 branch_block_stmt_13736/EQ_u1_u1_13959_place
      -- 
    e_block_daemon_CP_11105_elements(203) <= e_block_daemon_CP_11105_elements(202);
    -- CP-element group 204:  transition  bypass 
    -- CP-element group 204: predecessors 
    -- CP-element group 204: 	203 
    -- CP-element group 204: successors 
    -- CP-element group 204: 	205 
    -- CP-element group 204:  members (1) 
      -- CP-element group 204: 	 branch_block_stmt_13736/if_stmt_13956_if_link/$entry
      -- 
    e_block_daemon_CP_11105_elements(204) <= e_block_daemon_CP_11105_elements(203);
    -- CP-element group 205:  transition  input  bypass 
    -- CP-element group 205: predecessors 
    -- CP-element group 205: 	204 
    -- CP-element group 205: successors 
    -- CP-element group 205: 	208 
    -- CP-element group 205:  members (2) 
      -- CP-element group 205: 	 branch_block_stmt_13736/if_stmt_13956_if_link/if_choice_transition
      -- CP-element group 205: 	 branch_block_stmt_13736/if_stmt_13956_if_link/$exit
      -- 
    if_choice_transition_12194_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 205_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_13956_branch_ack_1, ack => e_block_daemon_CP_11105_elements(205)); -- 
    -- CP-element group 206:  transition  bypass 
    -- CP-element group 206: predecessors 
    -- CP-element group 206: 	203 
    -- CP-element group 206: successors 
    -- CP-element group 206: 	207 
    -- CP-element group 206:  members (1) 
      -- CP-element group 206: 	 branch_block_stmt_13736/if_stmt_13956_else_link/$entry
      -- 
    e_block_daemon_CP_11105_elements(206) <= e_block_daemon_CP_11105_elements(203);
    -- CP-element group 207:  transition  input  bypass 
    -- CP-element group 207: predecessors 
    -- CP-element group 207: 	206 
    -- CP-element group 207: successors 
    -- CP-element group 207: 	209 
    -- CP-element group 207:  members (2) 
      -- CP-element group 207: 	 branch_block_stmt_13736/if_stmt_13956_else_link/else_choice_transition
      -- CP-element group 207: 	 branch_block_stmt_13736/if_stmt_13956_else_link/$exit
      -- 
    else_choice_transition_12198_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 207_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_13956_branch_ack_0, ack => e_block_daemon_CP_11105_elements(207)); -- 
    -- CP-element group 208:  place  bypass 
    -- CP-element group 208: predecessors 
    -- CP-element group 208: 	205 
    -- CP-element group 208: successors 
    -- CP-element group 208: 	224 
    -- CP-element group 208:  members (1) 
      -- CP-element group 208: 	 branch_block_stmt_13736/GotNewKey
      -- 
    e_block_daemon_CP_11105_elements(208) <= e_block_daemon_CP_11105_elements(205);
    -- CP-element group 209:  place  bypass 
    -- CP-element group 209: predecessors 
    -- CP-element group 209: 	207 
    -- CP-element group 209: successors 
    -- CP-element group 209: 	242 
    -- CP-element group 209:  members (1) 
      -- CP-element group 209: 	 branch_block_stmt_13736/NotGotNewKey
      -- 
    e_block_daemon_CP_11105_elements(209) <= e_block_daemon_CP_11105_elements(207);
    -- CP-element group 210:  transition  bypass 
    -- CP-element group 210: predecessors 
    -- CP-element group 210: 	2 
    -- CP-element group 210: successors 
    -- CP-element group 210:  members (1) 
      -- CP-element group 210: 	 branch_block_stmt_13736/merge_stmt_13740_dead_link/$entry
      -- 
    e_block_daemon_CP_11105_elements(210) <= e_block_daemon_CP_11105_elements(2);
    -- CP-element group 211:  transition  bypass 
    -- CP-element group 211: predecessors 
    -- CP-element group 211: 	2 
    -- CP-element group 211: successors 
    -- CP-element group 211: 	213 
    -- CP-element group 211:  members (2) 
      -- CP-element group 211: 	 branch_block_stmt_13736/merge_stmt_13740__entry___PhiReq/$exit
      -- CP-element group 211: 	 branch_block_stmt_13736/merge_stmt_13740__entry___PhiReq/$entry
      -- 
    e_block_daemon_CP_11105_elements(211) <= e_block_daemon_CP_11105_elements(2);
    -- CP-element group 212:  transition  bypass 
    -- CP-element group 212: predecessors 
    -- CP-element group 212: 	28 
    -- CP-element group 212: successors 
    -- CP-element group 212: 	213 
    -- CP-element group 212:  members (2) 
      -- CP-element group 212: 	 branch_block_stmt_13736/NotGotCmd_PhiReq/$exit
      -- CP-element group 212: 	 branch_block_stmt_13736/NotGotCmd_PhiReq/$entry
      -- 
    e_block_daemon_CP_11105_elements(212) <= e_block_daemon_CP_11105_elements(28);
    -- CP-element group 213:  merge  place  bypass 
    -- CP-element group 213: predecessors 
    -- CP-element group 213: 	211 
    -- CP-element group 213: 	212 
    -- CP-element group 213: successors 
    -- CP-element group 213: 	214 
    -- CP-element group 213:  members (1) 
      -- CP-element group 213: 	 branch_block_stmt_13736/merge_stmt_13740_PhiReqMerge
      -- 
    e_block_daemon_CP_11105_elements(213) <= OrReduce(e_block_daemon_CP_11105_elements(211) & e_block_daemon_CP_11105_elements(212));
    -- CP-element group 214:  transition  bypass 
    -- CP-element group 214: predecessors 
    -- CP-element group 214: 	213 
    -- CP-element group 214: successors 
    -- CP-element group 214: 	3 
    -- CP-element group 214:  members (3) 
      -- CP-element group 214: 	 branch_block_stmt_13736/merge_stmt_13740_PhiAck/dummy
      -- CP-element group 214: 	 branch_block_stmt_13736/merge_stmt_13740_PhiAck/$exit
      -- CP-element group 214: 	 branch_block_stmt_13736/merge_stmt_13740_PhiAck/$entry
      -- 
    e_block_daemon_CP_11105_elements(214) <= e_block_daemon_CP_11105_elements(213);
    -- CP-element group 215:  transition  bypass 
    -- CP-element group 215: predecessors 
    -- CP-element group 215: 	6 
    -- CP-element group 215: successors 
    -- CP-element group 215:  members (1) 
      -- CP-element group 215: 	 branch_block_stmt_13736/merge_stmt_13762_dead_link/$entry
      -- 
    e_block_daemon_CP_11105_elements(215) <= e_block_daemon_CP_11105_elements(6);
    -- CP-element group 216:  fork  transition  output  bypass 
    -- CP-element group 216: predecessors 
    -- CP-element group 216: 	6 
    -- CP-element group 216: successors 
    -- CP-element group 216: 	217 
    -- CP-element group 216: 	218 
    -- CP-element group 216: 	220 
    -- CP-element group 216: 	221 
    -- CP-element group 216:  members (15) 
      -- CP-element group 216: 	 branch_block_stmt_13736/merge_stmt_13762__entry___PhiReq/phi_stmt_13767/phi_stmt_13767_sources/Interlock/$entry
      -- CP-element group 216: 	 branch_block_stmt_13736/merge_stmt_13762__entry___PhiReq/phi_stmt_13763/phi_stmt_13763_sources/Interlock/Update/req
      -- CP-element group 216: 	 branch_block_stmt_13736/merge_stmt_13762__entry___PhiReq/phi_stmt_13763/phi_stmt_13763_sources/Interlock/$entry
      -- CP-element group 216: 	 branch_block_stmt_13736/merge_stmt_13762__entry___PhiReq/phi_stmt_13767/phi_stmt_13767_sources/$entry
      -- CP-element group 216: 	 branch_block_stmt_13736/merge_stmt_13762__entry___PhiReq/phi_stmt_13767/$entry
      -- CP-element group 216: 	 branch_block_stmt_13736/merge_stmt_13762__entry___PhiReq/phi_stmt_13763/phi_stmt_13763_sources/Interlock/Sample/req
      -- CP-element group 216: 	 branch_block_stmt_13736/merge_stmt_13762__entry___PhiReq/phi_stmt_13767/phi_stmt_13767_sources/Interlock/Update/req
      -- CP-element group 216: 	 branch_block_stmt_13736/merge_stmt_13762__entry___PhiReq/phi_stmt_13763/phi_stmt_13763_sources/Interlock/Update/$entry
      -- CP-element group 216: 	 branch_block_stmt_13736/merge_stmt_13762__entry___PhiReq/phi_stmt_13767/phi_stmt_13767_sources/Interlock/Update/$entry
      -- CP-element group 216: 	 branch_block_stmt_13736/merge_stmt_13762__entry___PhiReq/phi_stmt_13763/phi_stmt_13763_sources/$entry
      -- CP-element group 216: 	 branch_block_stmt_13736/merge_stmt_13762__entry___PhiReq/phi_stmt_13763/$entry
      -- CP-element group 216: 	 branch_block_stmt_13736/merge_stmt_13762__entry___PhiReq/phi_stmt_13763/phi_stmt_13763_sources/Interlock/Sample/$entry
      -- CP-element group 216: 	 branch_block_stmt_13736/merge_stmt_13762__entry___PhiReq/$entry
      -- CP-element group 216: 	 branch_block_stmt_13736/merge_stmt_13762__entry___PhiReq/phi_stmt_13767/phi_stmt_13767_sources/Interlock/Sample/req
      -- CP-element group 216: 	 branch_block_stmt_13736/merge_stmt_13762__entry___PhiReq/phi_stmt_13767/phi_stmt_13767_sources/Interlock/Sample/$entry
      -- 
    req_12235_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_12235_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_block_daemon_CP_11105_elements(216), ack => e_init_key_13755_13765_buf_req_0); -- 
    req_12240_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_12240_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_block_daemon_CP_11105_elements(216), ack => e_init_key_13755_13765_buf_req_1); -- 
    req_12255_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_12255_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_block_daemon_CP_11105_elements(216), ack => e_init_count_13751_13769_buf_req_0); -- 
    req_12260_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_12260_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_block_daemon_CP_11105_elements(216), ack => e_init_count_13751_13769_buf_req_1); -- 
    e_block_daemon_CP_11105_elements(216) <= e_block_daemon_CP_11105_elements(6);
    -- CP-element group 217:  transition  input  bypass 
    -- CP-element group 217: predecessors 
    -- CP-element group 217: 	216 
    -- CP-element group 217: successors 
    -- CP-element group 217: 	219 
    -- CP-element group 217:  members (2) 
      -- CP-element group 217: 	 branch_block_stmt_13736/merge_stmt_13762__entry___PhiReq/phi_stmt_13763/phi_stmt_13763_sources/Interlock/Sample/ack
      -- CP-element group 217: 	 branch_block_stmt_13736/merge_stmt_13762__entry___PhiReq/phi_stmt_13763/phi_stmt_13763_sources/Interlock/Sample/$exit
      -- 
    ack_12236_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 217_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_init_key_13755_13765_buf_ack_0, ack => e_block_daemon_CP_11105_elements(217)); -- 
    -- CP-element group 218:  transition  input  bypass 
    -- CP-element group 218: predecessors 
    -- CP-element group 218: 	216 
    -- CP-element group 218: successors 
    -- CP-element group 218: 	219 
    -- CP-element group 218:  members (2) 
      -- CP-element group 218: 	 branch_block_stmt_13736/merge_stmt_13762__entry___PhiReq/phi_stmt_13763/phi_stmt_13763_sources/Interlock/Update/ack
      -- CP-element group 218: 	 branch_block_stmt_13736/merge_stmt_13762__entry___PhiReq/phi_stmt_13763/phi_stmt_13763_sources/Interlock/Update/$exit
      -- 
    ack_12241_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 218_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_init_key_13755_13765_buf_ack_1, ack => e_block_daemon_CP_11105_elements(218)); -- 
    -- CP-element group 219:  join  transition  output  bypass 
    -- CP-element group 219: predecessors 
    -- CP-element group 219: 	217 
    -- CP-element group 219: 	218 
    -- CP-element group 219: successors 
    -- CP-element group 219: 	223 
    -- CP-element group 219:  members (4) 
      -- CP-element group 219: 	 branch_block_stmt_13736/merge_stmt_13762__entry___PhiReq/phi_stmt_13763/phi_stmt_13763_sources/Interlock/$exit
      -- CP-element group 219: 	 branch_block_stmt_13736/merge_stmt_13762__entry___PhiReq/phi_stmt_13763/phi_stmt_13763_req
      -- CP-element group 219: 	 branch_block_stmt_13736/merge_stmt_13762__entry___PhiReq/phi_stmt_13763/phi_stmt_13763_sources/$exit
      -- CP-element group 219: 	 branch_block_stmt_13736/merge_stmt_13762__entry___PhiReq/phi_stmt_13763/$exit
      -- 
    phi_stmt_13763_req_12242_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_13763_req_12242_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_block_daemon_CP_11105_elements(219), ack => phi_stmt_13763_req_0); -- 
    e_block_daemon_cp_element_group_219: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "e_block_daemon_cp_element_group_219"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= e_block_daemon_CP_11105_elements(217) & e_block_daemon_CP_11105_elements(218);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => e_block_daemon_CP_11105_elements(219), clk => clk, reset => reset); --
    end block;
    -- CP-element group 220:  transition  input  bypass 
    -- CP-element group 220: predecessors 
    -- CP-element group 220: 	216 
    -- CP-element group 220: successors 
    -- CP-element group 220: 	222 
    -- CP-element group 220:  members (2) 
      -- CP-element group 220: 	 branch_block_stmt_13736/merge_stmt_13762__entry___PhiReq/phi_stmt_13767/phi_stmt_13767_sources/Interlock/Sample/ack
      -- CP-element group 220: 	 branch_block_stmt_13736/merge_stmt_13762__entry___PhiReq/phi_stmt_13767/phi_stmt_13767_sources/Interlock/Sample/$exit
      -- 
    ack_12256_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 220_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_init_count_13751_13769_buf_ack_0, ack => e_block_daemon_CP_11105_elements(220)); -- 
    -- CP-element group 221:  transition  input  bypass 
    -- CP-element group 221: predecessors 
    -- CP-element group 221: 	216 
    -- CP-element group 221: successors 
    -- CP-element group 221: 	222 
    -- CP-element group 221:  members (2) 
      -- CP-element group 221: 	 branch_block_stmt_13736/merge_stmt_13762__entry___PhiReq/phi_stmt_13767/phi_stmt_13767_sources/Interlock/Update/ack
      -- CP-element group 221: 	 branch_block_stmt_13736/merge_stmt_13762__entry___PhiReq/phi_stmt_13767/phi_stmt_13767_sources/Interlock/Update/$exit
      -- 
    ack_12261_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 221_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_init_count_13751_13769_buf_ack_1, ack => e_block_daemon_CP_11105_elements(221)); -- 
    -- CP-element group 222:  join  transition  output  bypass 
    -- CP-element group 222: predecessors 
    -- CP-element group 222: 	220 
    -- CP-element group 222: 	221 
    -- CP-element group 222: successors 
    -- CP-element group 222: 	223 
    -- CP-element group 222:  members (4) 
      -- CP-element group 222: 	 branch_block_stmt_13736/merge_stmt_13762__entry___PhiReq/phi_stmt_13767/phi_stmt_13767_sources/Interlock/$exit
      -- CP-element group 222: 	 branch_block_stmt_13736/merge_stmt_13762__entry___PhiReq/phi_stmt_13767/phi_stmt_13767_sources/$exit
      -- CP-element group 222: 	 branch_block_stmt_13736/merge_stmt_13762__entry___PhiReq/phi_stmt_13767/$exit
      -- CP-element group 222: 	 branch_block_stmt_13736/merge_stmt_13762__entry___PhiReq/phi_stmt_13767/phi_stmt_13767_req
      -- 
    phi_stmt_13767_req_12262_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_13767_req_12262_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_block_daemon_CP_11105_elements(222), ack => phi_stmt_13767_req_0); -- 
    e_block_daemon_cp_element_group_222: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "e_block_daemon_cp_element_group_222"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= e_block_daemon_CP_11105_elements(220) & e_block_daemon_CP_11105_elements(221);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => e_block_daemon_CP_11105_elements(222), clk => clk, reset => reset); --
    end block;
    -- CP-element group 223:  join  transition  bypass 
    -- CP-element group 223: predecessors 
    -- CP-element group 223: 	219 
    -- CP-element group 223: 	222 
    -- CP-element group 223: successors 
    -- CP-element group 223: 	232 
    -- CP-element group 223:  members (1) 
      -- CP-element group 223: 	 branch_block_stmt_13736/merge_stmt_13762__entry___PhiReq/$exit
      -- 
    e_block_daemon_cp_element_group_223: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "e_block_daemon_cp_element_group_223"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= e_block_daemon_CP_11105_elements(219) & e_block_daemon_CP_11105_elements(222);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => e_block_daemon_CP_11105_elements(223), clk => clk, reset => reset); --
    end block;
    -- CP-element group 224:  fork  transition  output  bypass 
    -- CP-element group 224: predecessors 
    -- CP-element group 224: 	208 
    -- CP-element group 224: successors 
    -- CP-element group 224: 	225 
    -- CP-element group 224: 	226 
    -- CP-element group 224: 	228 
    -- CP-element group 224: 	229 
    -- CP-element group 224:  members (15) 
      -- CP-element group 224: 	 branch_block_stmt_13736/GotNewKey_PhiReq/phi_stmt_13763/phi_stmt_13763_sources/Interlock/Update/req
      -- CP-element group 224: 	 branch_block_stmt_13736/GotNewKey_PhiReq/phi_stmt_13763/phi_stmt_13763_sources/Interlock/Update/$entry
      -- CP-element group 224: 	 branch_block_stmt_13736/GotNewKey_PhiReq/phi_stmt_13763/$entry
      -- CP-element group 224: 	 branch_block_stmt_13736/GotNewKey_PhiReq/$entry
      -- CP-element group 224: 	 branch_block_stmt_13736/GotNewKey_PhiReq/phi_stmt_13763/phi_stmt_13763_sources/Interlock/Sample/req
      -- CP-element group 224: 	 branch_block_stmt_13736/GotNewKey_PhiReq/phi_stmt_13767/phi_stmt_13767_sources/Interlock/Sample/req
      -- CP-element group 224: 	 branch_block_stmt_13736/GotNewKey_PhiReq/phi_stmt_13767/phi_stmt_13767_sources/Interlock/Sample/$entry
      -- CP-element group 224: 	 branch_block_stmt_13736/GotNewKey_PhiReq/phi_stmt_13763/phi_stmt_13763_sources/Interlock/Sample/$entry
      -- CP-element group 224: 	 branch_block_stmt_13736/GotNewKey_PhiReq/phi_stmt_13763/phi_stmt_13763_sources/Interlock/$entry
      -- CP-element group 224: 	 branch_block_stmt_13736/GotNewKey_PhiReq/phi_stmt_13767/phi_stmt_13767_sources/Interlock/$entry
      -- CP-element group 224: 	 branch_block_stmt_13736/GotNewKey_PhiReq/phi_stmt_13767/phi_stmt_13767_sources/$entry
      -- CP-element group 224: 	 branch_block_stmt_13736/GotNewKey_PhiReq/phi_stmt_13763/phi_stmt_13763_sources/$entry
      -- CP-element group 224: 	 branch_block_stmt_13736/GotNewKey_PhiReq/phi_stmt_13767/$entry
      -- CP-element group 224: 	 branch_block_stmt_13736/GotNewKey_PhiReq/phi_stmt_13767/phi_stmt_13767_sources/Interlock/Update/req
      -- CP-element group 224: 	 branch_block_stmt_13736/GotNewKey_PhiReq/phi_stmt_13767/phi_stmt_13767_sources/Interlock/Update/$entry
      -- 
    req_12278_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_12278_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_block_daemon_CP_11105_elements(224), ack => e_new_key_13955_13766_buf_req_0); -- 
    req_12283_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_12283_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_block_daemon_CP_11105_elements(224), ack => e_new_key_13955_13766_buf_req_1); -- 
    req_12298_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_12298_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_block_daemon_CP_11105_elements(224), ack => e_new_count_13951_13770_buf_req_0); -- 
    req_12303_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_12303_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_block_daemon_CP_11105_elements(224), ack => e_new_count_13951_13770_buf_req_1); -- 
    e_block_daemon_CP_11105_elements(224) <= e_block_daemon_CP_11105_elements(208);
    -- CP-element group 225:  transition  input  bypass 
    -- CP-element group 225: predecessors 
    -- CP-element group 225: 	224 
    -- CP-element group 225: successors 
    -- CP-element group 225: 	227 
    -- CP-element group 225:  members (2) 
      -- CP-element group 225: 	 branch_block_stmt_13736/GotNewKey_PhiReq/phi_stmt_13763/phi_stmt_13763_sources/Interlock/Sample/ack
      -- CP-element group 225: 	 branch_block_stmt_13736/GotNewKey_PhiReq/phi_stmt_13763/phi_stmt_13763_sources/Interlock/Sample/$exit
      -- 
    ack_12279_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 225_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_new_key_13955_13766_buf_ack_0, ack => e_block_daemon_CP_11105_elements(225)); -- 
    -- CP-element group 226:  transition  input  bypass 
    -- CP-element group 226: predecessors 
    -- CP-element group 226: 	224 
    -- CP-element group 226: successors 
    -- CP-element group 226: 	227 
    -- CP-element group 226:  members (2) 
      -- CP-element group 226: 	 branch_block_stmt_13736/GotNewKey_PhiReq/phi_stmt_13763/phi_stmt_13763_sources/Interlock/Update/$exit
      -- CP-element group 226: 	 branch_block_stmt_13736/GotNewKey_PhiReq/phi_stmt_13763/phi_stmt_13763_sources/Interlock/Update/ack
      -- 
    ack_12284_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 226_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_new_key_13955_13766_buf_ack_1, ack => e_block_daemon_CP_11105_elements(226)); -- 
    -- CP-element group 227:  join  transition  output  bypass 
    -- CP-element group 227: predecessors 
    -- CP-element group 227: 	225 
    -- CP-element group 227: 	226 
    -- CP-element group 227: successors 
    -- CP-element group 227: 	231 
    -- CP-element group 227:  members (4) 
      -- CP-element group 227: 	 branch_block_stmt_13736/GotNewKey_PhiReq/phi_stmt_13763/phi_stmt_13763_sources/Interlock/$exit
      -- CP-element group 227: 	 branch_block_stmt_13736/GotNewKey_PhiReq/phi_stmt_13763/phi_stmt_13763_sources/$exit
      -- CP-element group 227: 	 branch_block_stmt_13736/GotNewKey_PhiReq/phi_stmt_13763/phi_stmt_13763_req
      -- CP-element group 227: 	 branch_block_stmt_13736/GotNewKey_PhiReq/phi_stmt_13763/$exit
      -- 
    phi_stmt_13763_req_12285_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_13763_req_12285_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_block_daemon_CP_11105_elements(227), ack => phi_stmt_13763_req_1); -- 
    e_block_daemon_cp_element_group_227: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "e_block_daemon_cp_element_group_227"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= e_block_daemon_CP_11105_elements(225) & e_block_daemon_CP_11105_elements(226);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => e_block_daemon_CP_11105_elements(227), clk => clk, reset => reset); --
    end block;
    -- CP-element group 228:  transition  input  bypass 
    -- CP-element group 228: predecessors 
    -- CP-element group 228: 	224 
    -- CP-element group 228: successors 
    -- CP-element group 228: 	230 
    -- CP-element group 228:  members (2) 
      -- CP-element group 228: 	 branch_block_stmt_13736/GotNewKey_PhiReq/phi_stmt_13767/phi_stmt_13767_sources/Interlock/Sample/ack
      -- CP-element group 228: 	 branch_block_stmt_13736/GotNewKey_PhiReq/phi_stmt_13767/phi_stmt_13767_sources/Interlock/Sample/$exit
      -- 
    ack_12299_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 228_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_new_count_13951_13770_buf_ack_0, ack => e_block_daemon_CP_11105_elements(228)); -- 
    -- CP-element group 229:  transition  input  bypass 
    -- CP-element group 229: predecessors 
    -- CP-element group 229: 	224 
    -- CP-element group 229: successors 
    -- CP-element group 229: 	230 
    -- CP-element group 229:  members (2) 
      -- CP-element group 229: 	 branch_block_stmt_13736/GotNewKey_PhiReq/phi_stmt_13767/phi_stmt_13767_sources/Interlock/Update/ack
      -- CP-element group 229: 	 branch_block_stmt_13736/GotNewKey_PhiReq/phi_stmt_13767/phi_stmt_13767_sources/Interlock/Update/$exit
      -- 
    ack_12304_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 229_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_new_count_13951_13770_buf_ack_1, ack => e_block_daemon_CP_11105_elements(229)); -- 
    -- CP-element group 230:  join  transition  output  bypass 
    -- CP-element group 230: predecessors 
    -- CP-element group 230: 	228 
    -- CP-element group 230: 	229 
    -- CP-element group 230: successors 
    -- CP-element group 230: 	231 
    -- CP-element group 230:  members (4) 
      -- CP-element group 230: 	 branch_block_stmt_13736/GotNewKey_PhiReq/phi_stmt_13767/phi_stmt_13767_sources/Interlock/$exit
      -- CP-element group 230: 	 branch_block_stmt_13736/GotNewKey_PhiReq/phi_stmt_13767/phi_stmt_13767_req
      -- CP-element group 230: 	 branch_block_stmt_13736/GotNewKey_PhiReq/phi_stmt_13767/phi_stmt_13767_sources/$exit
      -- CP-element group 230: 	 branch_block_stmt_13736/GotNewKey_PhiReq/phi_stmt_13767/$exit
      -- 
    phi_stmt_13767_req_12305_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_13767_req_12305_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_block_daemon_CP_11105_elements(230), ack => phi_stmt_13767_req_1); -- 
    e_block_daemon_cp_element_group_230: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "e_block_daemon_cp_element_group_230"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= e_block_daemon_CP_11105_elements(228) & e_block_daemon_CP_11105_elements(229);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => e_block_daemon_CP_11105_elements(230), clk => clk, reset => reset); --
    end block;
    -- CP-element group 231:  join  transition  bypass 
    -- CP-element group 231: predecessors 
    -- CP-element group 231: 	227 
    -- CP-element group 231: 	230 
    -- CP-element group 231: successors 
    -- CP-element group 231: 	232 
    -- CP-element group 231:  members (1) 
      -- CP-element group 231: 	 branch_block_stmt_13736/GotNewKey_PhiReq/$exit
      -- 
    e_block_daemon_cp_element_group_231: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "e_block_daemon_cp_element_group_231"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= e_block_daemon_CP_11105_elements(227) & e_block_daemon_CP_11105_elements(230);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => e_block_daemon_CP_11105_elements(231), clk => clk, reset => reset); --
    end block;
    -- CP-element group 232:  merge  place  bypass 
    -- CP-element group 232: predecessors 
    -- CP-element group 232: 	223 
    -- CP-element group 232: 	231 
    -- CP-element group 232: successors 
    -- CP-element group 232: 	233 
    -- CP-element group 232:  members (1) 
      -- CP-element group 232: 	 branch_block_stmt_13736/merge_stmt_13762_PhiReqMerge
      -- 
    e_block_daemon_CP_11105_elements(232) <= OrReduce(e_block_daemon_CP_11105_elements(223) & e_block_daemon_CP_11105_elements(231));
    -- CP-element group 233:  fork  transition  bypass 
    -- CP-element group 233: predecessors 
    -- CP-element group 233: 	232 
    -- CP-element group 233: successors 
    -- CP-element group 233: 	234 
    -- CP-element group 233: 	235 
    -- CP-element group 233:  members (1) 
      -- CP-element group 233: 	 branch_block_stmt_13736/merge_stmt_13762_PhiAck/$entry
      -- 
    e_block_daemon_CP_11105_elements(233) <= e_block_daemon_CP_11105_elements(232);
    -- CP-element group 234:  transition  input  bypass 
    -- CP-element group 234: predecessors 
    -- CP-element group 234: 	233 
    -- CP-element group 234: successors 
    -- CP-element group 234: 	236 
    -- CP-element group 234:  members (1) 
      -- CP-element group 234: 	 branch_block_stmt_13736/merge_stmt_13762_PhiAck/phi_stmt_13763_ack
      -- 
    phi_stmt_13763_ack_12310_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 234_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_13763_ack_0, ack => e_block_daemon_CP_11105_elements(234)); -- 
    -- CP-element group 235:  transition  input  bypass 
    -- CP-element group 235: predecessors 
    -- CP-element group 235: 	233 
    -- CP-element group 235: successors 
    -- CP-element group 235: 	236 
    -- CP-element group 235:  members (1) 
      -- CP-element group 235: 	 branch_block_stmt_13736/merge_stmt_13762_PhiAck/phi_stmt_13767_ack
      -- 
    phi_stmt_13767_ack_12311_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 235_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_13767_ack_0, ack => e_block_daemon_CP_11105_elements(235)); -- 
    -- CP-element group 236:  join  transition  bypass 
    -- CP-element group 236: predecessors 
    -- CP-element group 236: 	234 
    -- CP-element group 236: 	235 
    -- CP-element group 236: successors 
    -- CP-element group 236: 	7 
    -- CP-element group 236:  members (1) 
      -- CP-element group 236: 	 branch_block_stmt_13736/merge_stmt_13762_PhiAck/$exit
      -- 
    e_block_daemon_cp_element_group_236: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "e_block_daemon_cp_element_group_236"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= e_block_daemon_CP_11105_elements(234) & e_block_daemon_CP_11105_elements(235);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => e_block_daemon_CP_11105_elements(236), clk => clk, reset => reset); --
    end block;
    -- CP-element group 237:  transition  bypass 
    -- CP-element group 237: predecessors 
    -- CP-element group 237: 	8 
    -- CP-element group 237: successors 
    -- CP-element group 237:  members (1) 
      -- CP-element group 237: 	 branch_block_stmt_13736/merge_stmt_13822_dead_link/$entry
      -- 
    e_block_daemon_CP_11105_elements(237) <= e_block_daemon_CP_11105_elements(8);
    -- CP-element group 238:  fork  transition  output  bypass 
    -- CP-element group 238: predecessors 
    -- CP-element group 238: 	8 
    -- CP-element group 238: successors 
    -- CP-element group 238: 	239 
    -- CP-element group 238: 	240 
    -- CP-element group 238:  members (8) 
      -- CP-element group 238: 	 branch_block_stmt_13736/merge_stmt_13822__entry___PhiReq/phi_stmt_13823/phi_stmt_13823_sources/$entry
      -- CP-element group 238: 	 branch_block_stmt_13736/merge_stmt_13822__entry___PhiReq/phi_stmt_13823/phi_stmt_13823_sources/Interlock/$entry
      -- CP-element group 238: 	 branch_block_stmt_13736/merge_stmt_13822__entry___PhiReq/phi_stmt_13823/$entry
      -- CP-element group 238: 	 branch_block_stmt_13736/merge_stmt_13822__entry___PhiReq/phi_stmt_13823/phi_stmt_13823_sources/Interlock/Sample/$entry
      -- CP-element group 238: 	 branch_block_stmt_13736/merge_stmt_13822__entry___PhiReq/$entry
      -- CP-element group 238: 	 branch_block_stmt_13736/merge_stmt_13822__entry___PhiReq/phi_stmt_13823/phi_stmt_13823_sources/Interlock/Sample/req
      -- CP-element group 238: 	 branch_block_stmt_13736/merge_stmt_13822__entry___PhiReq/phi_stmt_13823/phi_stmt_13823_sources/Interlock/Update/$entry
      -- CP-element group 238: 	 branch_block_stmt_13736/merge_stmt_13822__entry___PhiReq/phi_stmt_13823/phi_stmt_13823_sources/Interlock/Update/req
      -- 
    req_12331_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_12331_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_block_daemon_CP_11105_elements(238), ack => countA_13767_13825_buf_req_0); -- 
    req_12336_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_12336_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_block_daemon_CP_11105_elements(238), ack => countA_13767_13825_buf_req_1); -- 
    e_block_daemon_CP_11105_elements(238) <= e_block_daemon_CP_11105_elements(8);
    -- CP-element group 239:  transition  input  bypass 
    -- CP-element group 239: predecessors 
    -- CP-element group 239: 	238 
    -- CP-element group 239: successors 
    -- CP-element group 239: 	241 
    -- CP-element group 239:  members (2) 
      -- CP-element group 239: 	 branch_block_stmt_13736/merge_stmt_13822__entry___PhiReq/phi_stmt_13823/phi_stmt_13823_sources/Interlock/Sample/$exit
      -- CP-element group 239: 	 branch_block_stmt_13736/merge_stmt_13822__entry___PhiReq/phi_stmt_13823/phi_stmt_13823_sources/Interlock/Sample/ack
      -- 
    ack_12332_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 239_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => countA_13767_13825_buf_ack_0, ack => e_block_daemon_CP_11105_elements(239)); -- 
    -- CP-element group 240:  transition  input  bypass 
    -- CP-element group 240: predecessors 
    -- CP-element group 240: 	238 
    -- CP-element group 240: successors 
    -- CP-element group 240: 	241 
    -- CP-element group 240:  members (2) 
      -- CP-element group 240: 	 branch_block_stmt_13736/merge_stmt_13822__entry___PhiReq/phi_stmt_13823/phi_stmt_13823_sources/Interlock/Update/$exit
      -- CP-element group 240: 	 branch_block_stmt_13736/merge_stmt_13822__entry___PhiReq/phi_stmt_13823/phi_stmt_13823_sources/Interlock/Update/ack
      -- 
    ack_12337_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 240_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => countA_13767_13825_buf_ack_1, ack => e_block_daemon_CP_11105_elements(240)); -- 
    -- CP-element group 241:  join  transition  output  bypass 
    -- CP-element group 241: predecessors 
    -- CP-element group 241: 	239 
    -- CP-element group 241: 	240 
    -- CP-element group 241: successors 
    -- CP-element group 241: 	246 
    -- CP-element group 241:  members (5) 
      -- CP-element group 241: 	 branch_block_stmt_13736/merge_stmt_13822__entry___PhiReq/phi_stmt_13823/phi_stmt_13823_sources/$exit
      -- CP-element group 241: 	 branch_block_stmt_13736/merge_stmt_13822__entry___PhiReq/phi_stmt_13823/phi_stmt_13823_sources/Interlock/$exit
      -- CP-element group 241: 	 branch_block_stmt_13736/merge_stmt_13822__entry___PhiReq/phi_stmt_13823/$exit
      -- CP-element group 241: 	 branch_block_stmt_13736/merge_stmt_13822__entry___PhiReq/$exit
      -- CP-element group 241: 	 branch_block_stmt_13736/merge_stmt_13822__entry___PhiReq/phi_stmt_13823/phi_stmt_13823_req
      -- 
    phi_stmt_13823_req_12338_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_13823_req_12338_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_block_daemon_CP_11105_elements(241), ack => phi_stmt_13823_req_0); -- 
    e_block_daemon_cp_element_group_241: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "e_block_daemon_cp_element_group_241"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= e_block_daemon_CP_11105_elements(239) & e_block_daemon_CP_11105_elements(240);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => e_block_daemon_CP_11105_elements(241), clk => clk, reset => reset); --
    end block;
    -- CP-element group 242:  fork  transition  output  bypass 
    -- CP-element group 242: predecessors 
    -- CP-element group 242: 	209 
    -- CP-element group 242: successors 
    -- CP-element group 242: 	243 
    -- CP-element group 242: 	244 
    -- CP-element group 242:  members (8) 
      -- CP-element group 242: 	 branch_block_stmt_13736/NotGotNewKey_PhiReq/$entry
      -- CP-element group 242: 	 branch_block_stmt_13736/NotGotNewKey_PhiReq/phi_stmt_13823/$entry
      -- CP-element group 242: 	 branch_block_stmt_13736/NotGotNewKey_PhiReq/phi_stmt_13823/phi_stmt_13823_sources/$entry
      -- CP-element group 242: 	 branch_block_stmt_13736/NotGotNewKey_PhiReq/phi_stmt_13823/phi_stmt_13823_sources/Interlock/$entry
      -- CP-element group 242: 	 branch_block_stmt_13736/NotGotNewKey_PhiReq/phi_stmt_13823/phi_stmt_13823_sources/Interlock/Sample/$entry
      -- CP-element group 242: 	 branch_block_stmt_13736/NotGotNewKey_PhiReq/phi_stmt_13823/phi_stmt_13823_sources/Interlock/Sample/req
      -- CP-element group 242: 	 branch_block_stmt_13736/NotGotNewKey_PhiReq/phi_stmt_13823/phi_stmt_13823_sources/Interlock/Update/$entry
      -- CP-element group 242: 	 branch_block_stmt_13736/NotGotNewKey_PhiReq/phi_stmt_13823/phi_stmt_13823_sources/Interlock/Update/req
      -- 
    req_12354_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_12354_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_block_daemon_CP_11105_elements(242), ack => e_new_count_13951_13826_buf_req_0); -- 
    req_12359_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_12359_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_block_daemon_CP_11105_elements(242), ack => e_new_count_13951_13826_buf_req_1); -- 
    e_block_daemon_CP_11105_elements(242) <= e_block_daemon_CP_11105_elements(209);
    -- CP-element group 243:  transition  input  bypass 
    -- CP-element group 243: predecessors 
    -- CP-element group 243: 	242 
    -- CP-element group 243: successors 
    -- CP-element group 243: 	245 
    -- CP-element group 243:  members (2) 
      -- CP-element group 243: 	 branch_block_stmt_13736/NotGotNewKey_PhiReq/phi_stmt_13823/phi_stmt_13823_sources/Interlock/Sample/$exit
      -- CP-element group 243: 	 branch_block_stmt_13736/NotGotNewKey_PhiReq/phi_stmt_13823/phi_stmt_13823_sources/Interlock/Sample/ack
      -- 
    ack_12355_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 243_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_new_count_13951_13826_buf_ack_0, ack => e_block_daemon_CP_11105_elements(243)); -- 
    -- CP-element group 244:  transition  input  bypass 
    -- CP-element group 244: predecessors 
    -- CP-element group 244: 	242 
    -- CP-element group 244: successors 
    -- CP-element group 244: 	245 
    -- CP-element group 244:  members (2) 
      -- CP-element group 244: 	 branch_block_stmt_13736/NotGotNewKey_PhiReq/phi_stmt_13823/phi_stmt_13823_sources/Interlock/Update/$exit
      -- CP-element group 244: 	 branch_block_stmt_13736/NotGotNewKey_PhiReq/phi_stmt_13823/phi_stmt_13823_sources/Interlock/Update/ack
      -- 
    ack_12360_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 244_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_new_count_13951_13826_buf_ack_1, ack => e_block_daemon_CP_11105_elements(244)); -- 
    -- CP-element group 245:  join  transition  output  bypass 
    -- CP-element group 245: predecessors 
    -- CP-element group 245: 	243 
    -- CP-element group 245: 	244 
    -- CP-element group 245: successors 
    -- CP-element group 245: 	246 
    -- CP-element group 245:  members (5) 
      -- CP-element group 245: 	 branch_block_stmt_13736/NotGotNewKey_PhiReq/$exit
      -- CP-element group 245: 	 branch_block_stmt_13736/NotGotNewKey_PhiReq/phi_stmt_13823/$exit
      -- CP-element group 245: 	 branch_block_stmt_13736/NotGotNewKey_PhiReq/phi_stmt_13823/phi_stmt_13823_sources/$exit
      -- CP-element group 245: 	 branch_block_stmt_13736/NotGotNewKey_PhiReq/phi_stmt_13823/phi_stmt_13823_sources/Interlock/$exit
      -- CP-element group 245: 	 branch_block_stmt_13736/NotGotNewKey_PhiReq/phi_stmt_13823/phi_stmt_13823_req
      -- 
    phi_stmt_13823_req_12361_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_13823_req_12361_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => e_block_daemon_CP_11105_elements(245), ack => phi_stmt_13823_req_1); -- 
    e_block_daemon_cp_element_group_245: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "e_block_daemon_cp_element_group_245"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= e_block_daemon_CP_11105_elements(243) & e_block_daemon_CP_11105_elements(244);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => e_block_daemon_CP_11105_elements(245), clk => clk, reset => reset); --
    end block;
    -- CP-element group 246:  merge  place  bypass 
    -- CP-element group 246: predecessors 
    -- CP-element group 246: 	241 
    -- CP-element group 246: 	245 
    -- CP-element group 246: successors 
    -- CP-element group 246: 	247 
    -- CP-element group 246:  members (1) 
      -- CP-element group 246: 	 branch_block_stmt_13736/merge_stmt_13822_PhiReqMerge
      -- 
    e_block_daemon_CP_11105_elements(246) <= OrReduce(e_block_daemon_CP_11105_elements(241) & e_block_daemon_CP_11105_elements(245));
    -- CP-element group 247:  transition  bypass 
    -- CP-element group 247: predecessors 
    -- CP-element group 247: 	246 
    -- CP-element group 247: successors 
    -- CP-element group 247: 	248 
    -- CP-element group 247:  members (1) 
      -- CP-element group 247: 	 branch_block_stmt_13736/merge_stmt_13822_PhiAck/$entry
      -- 
    e_block_daemon_CP_11105_elements(247) <= e_block_daemon_CP_11105_elements(246);
    -- CP-element group 248:  transition  input  bypass 
    -- CP-element group 248: predecessors 
    -- CP-element group 248: 	247 
    -- CP-element group 248: successors 
    -- CP-element group 248: 	9 
    -- CP-element group 248:  members (2) 
      -- CP-element group 248: 	 branch_block_stmt_13736/merge_stmt_13822_PhiAck/$exit
      -- CP-element group 248: 	 branch_block_stmt_13736/merge_stmt_13822_PhiAck/phi_stmt_13823_ack
      -- 
    phi_stmt_13823_ack_12366_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 248_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_13823_ack_0, ack => e_block_daemon_CP_11105_elements(248)); -- 
    -- CP-element group 249:  join  transition  bypass  pipeline-parent 
    -- CP-element group 249: predecessors 
    -- CP-element group 249: 	183 
    -- CP-element group 249: 	71 
    -- CP-element group 249: successors 
    -- CP-element group 249: 	55 
    -- CP-element group 249:  members (2) 
      -- CP-element group 249: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/$exit
      -- CP-element group 249: 	 branch_block_stmt_13736/do_while_stmt_13828/do_while_stmt_13828_loop_body/phi_stmt_13830_phi_mux_ack_ps
      -- 
    e_block_daemon_cp_element_group_249: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 2,1 => 2);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "e_block_daemon_cp_element_group_249"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= e_block_daemon_CP_11105_elements(183) & e_block_daemon_CP_11105_elements(71);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => e_block_daemon_CP_11105_elements(249), clk => clk, reset => reset); --
    end block;
    do_while_stmt_13828_terminator_12071: loop_terminator -- 
      generic map (name => " do_while_stmt_13828_terminator_12071", max_iterations_in_flight =>2) 
      port map(loop_body_exit => e_block_daemon_CP_11105_elements(55),loop_continue => e_block_daemon_CP_11105_elements(192),loop_terminate => e_block_daemon_CP_11105_elements(190),loop_back => e_block_daemon_CP_11105_elements(53),loop_exit => e_block_daemon_CP_11105_elements(52),clk => clk, reset => reset); -- 
    phi_stmt_13830_phi_seq_11550_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= e_block_daemon_CP_11105_elements(66);
      e_block_daemon_CP_11105_elements(72)<= src_sample_reqs(0);
      src_sample_acks(0)  <= e_block_daemon_CP_11105_elements(72);
      e_block_daemon_CP_11105_elements(73)<= src_update_reqs(0);
      src_update_acks(0)  <= e_block_daemon_CP_11105_elements(74);
      e_block_daemon_CP_11105_elements(67) <= phi_mux_reqs(0);
      triggers(1)  <= e_block_daemon_CP_11105_elements(64);
      e_block_daemon_CP_11105_elements(76)<= src_sample_reqs(1);
      src_sample_acks(1)  <= e_block_daemon_CP_11105_elements(78);
      e_block_daemon_CP_11105_elements(77)<= src_update_reqs(1);
      src_update_acks(1)  <= e_block_daemon_CP_11105_elements(79);
      e_block_daemon_CP_11105_elements(65) <= phi_mux_reqs(1);
      phi_stmt_13830_phi_seq_11550 : phi_sequencer_v2-- 
        generic map (place_capacity => 2, ntriggers => 2, name => "phi_stmt_13830_phi_seq_11550") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => e_block_daemon_CP_11105_elements(60), 
          phi_sample_ack => e_block_daemon_CP_11105_elements(62), 
          phi_update_req => e_block_daemon_CP_11105_elements(61), 
          phi_update_ack => e_block_daemon_CP_11105_elements(63), 
          phi_mux_ack => e_block_daemon_CP_11105_elements(71), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_11501_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= e_block_daemon_CP_11105_elements(56);
        preds(1)  <= e_block_daemon_CP_11105_elements(57);
        entry_tmerge_11501 : transition_merge -- 
          generic map(name => " entry_tmerge_11501")
          port map (preds => preds, symbol_out => e_block_daemon_CP_11105_elements(58));
          -- 
    end block;
    phi_stmt_13830_req_merge_11521_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= e_block_daemon_CP_11105_elements(69);
        preds(1)  <= e_block_daemon_CP_11105_elements(70);
        phi_stmt_13830_req_merge_11521 : transition_merge -- 
          generic map(name => " phi_stmt_13830_req_merge_11521")
          port map (preds => preds, symbol_out => e_block_daemon_CP_11105_elements(68));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal EQ_u1_u1_13759_wire : std_logic_vector(0 downto 0);
    signal EQ_u1_u1_13959_wire : std_logic_vector(0 downto 0);
    signal K0_13763 : std_logic_vector(127 downto 0);
    signal K10_13821 : std_logic_vector(127 downto 0);
    signal K10_13856_delayed_10_13920 : std_logic_vector(127 downto 0);
    signal K1_13776 : std_logic_vector(127 downto 0);
    signal K1_13811_delayed_1_13848 : std_logic_vector(127 downto 0);
    signal K2_13781 : std_logic_vector(127 downto 0);
    signal K2_13816_delayed_2_13856 : std_logic_vector(127 downto 0);
    signal K3_13786 : std_logic_vector(127 downto 0);
    signal K3_13821_delayed_3_13864 : std_logic_vector(127 downto 0);
    signal K4_13791 : std_logic_vector(127 downto 0);
    signal K4_13826_delayed_4_13872 : std_logic_vector(127 downto 0);
    signal K5_13796 : std_logic_vector(127 downto 0);
    signal K5_13831_delayed_5_13880 : std_logic_vector(127 downto 0);
    signal K6_13801 : std_logic_vector(127 downto 0);
    signal K6_13836_delayed_6_13888 : std_logic_vector(127 downto 0);
    signal K7_13806 : std_logic_vector(127 downto 0);
    signal K7_13841_delayed_7_13896 : std_logic_vector(127 downto 0);
    signal K8_13811 : std_logic_vector(127 downto 0);
    signal K8_13846_delayed_8_13904 : std_logic_vector(127 downto 0);
    signal K9_13816 : std_logic_vector(127 downto 0);
    signal K9_13851_delayed_9_13912 : std_logic_vector(127 downto 0);
    signal RConstant_10_13816 : std_logic_vector(7 downto 0);
    signal RConstant_11_13821 : std_logic_vector(7 downto 0);
    signal RConstant_2_13776 : std_logic_vector(7 downto 0);
    signal RConstant_3_13781 : std_logic_vector(7 downto 0);
    signal RConstant_4_13786 : std_logic_vector(7 downto 0);
    signal RConstant_5_13791 : std_logic_vector(7 downto 0);
    signal RConstant_6_13796 : std_logic_vector(7 downto 0);
    signal RConstant_7_13801 : std_logic_vector(7 downto 0);
    signal RConstant_8_13806 : std_logic_vector(7 downto 0);
    signal RConstant_9_13811 : std_logic_vector(7 downto 0);
    signal R_LAST_13923_wire_constant : std_logic_vector(0 downto 0);
    signal R_NOT_LAST_13851_wire_constant : std_logic_vector(0 downto 0);
    signal R_NOT_LAST_13859_wire_constant : std_logic_vector(0 downto 0);
    signal R_NOT_LAST_13867_wire_constant : std_logic_vector(0 downto 0);
    signal R_NOT_LAST_13875_wire_constant : std_logic_vector(0 downto 0);
    signal R_NOT_LAST_13883_wire_constant : std_logic_vector(0 downto 0);
    signal R_NOT_LAST_13891_wire_constant : std_logic_vector(0 downto 0);
    signal R_NOT_LAST_13899_wire_constant : std_logic_vector(0 downto 0);
    signal R_NOT_LAST_13907_wire_constant : std_logic_vector(0 downto 0);
    signal R_NOT_LAST_13915_wire_constant : std_logic_vector(0 downto 0);
    signal R_RConstant_1_13773_wire_constant : std_logic_vector(7 downto 0);
    signal R_ZERO_COUNT_13832_wire_constant : std_logic_vector(14 downto 0);
    signal ULT_u15_u1_13937_wire : std_logic_vector(0 downto 0);
    signal countA_13767 : std_logic_vector(14 downto 0);
    signal countA_13767_13825_buffered : std_logic_vector(14 downto 0);
    signal countB_13823 : std_logic_vector(14 downto 0);
    signal count_var_13830 : std_logic_vector(14 downto 0);
    signal e_get_key_13747 : std_logic_vector(0 downto 0);
    signal e_get_new_key_13947 : std_logic_vector(0 downto 0);
    signal e_init_cmd_13743 : std_logic_vector(143 downto 0);
    signal e_init_count_13751 : std_logic_vector(14 downto 0);
    signal e_init_count_13751_13769_buffered : std_logic_vector(14 downto 0);
    signal e_init_key_13755 : std_logic_vector(127 downto 0);
    signal e_init_key_13755_13765_buffered : std_logic_vector(127 downto 0);
    signal e_new_cmd_13943 : std_logic_vector(143 downto 0);
    signal e_new_count_13951 : std_logic_vector(14 downto 0);
    signal e_new_count_13951_13770_buffered : std_logic_vector(14 downto 0);
    signal e_new_count_13951_13826_buffered : std_logic_vector(14 downto 0);
    signal e_new_key_13955 : std_logic_vector(127 downto 0);
    signal e_new_key_13955_13766_buffered : std_logic_vector(127 downto 0);
    signal in128_13837 : std_logic_vector(127 downto 0);
    signal konst_13738_wire_constant : std_logic_vector(0 downto 0);
    signal konst_13758_wire_constant : std_logic_vector(0 downto 0);
    signal konst_13931_wire_constant : std_logic_vector(14 downto 0);
    signal konst_13939_wire_constant : std_logic_vector(0 downto 0);
    signal konst_13958_wire_constant : std_logic_vector(0 downto 0);
    signal n_count_var_13933 : std_logic_vector(14 downto 0);
    signal n_count_var_13933_13833_buffered : std_logic_vector(14 downto 0);
    signal round_S0_13810_delayed_1_13845 : std_logic_vector(127 downto 0);
    signal round_S0_13842 : std_logic_vector(127 downto 0);
    signal round_S10_13925 : std_logic_vector(127 downto 0);
    signal round_S1_13853 : std_logic_vector(127 downto 0);
    signal round_S2_13861 : std_logic_vector(127 downto 0);
    signal round_S3_13869 : std_logic_vector(127 downto 0);
    signal round_S4_13877 : std_logic_vector(127 downto 0);
    signal round_S5_13885 : std_logic_vector(127 downto 0);
    signal round_S6_13893 : std_logic_vector(127 downto 0);
    signal round_S7_13901 : std_logic_vector(127 downto 0);
    signal round_S8_13909 : std_logic_vector(127 downto 0);
    signal round_S9_13917 : std_logic_vector(127 downto 0);
    signal xxe_block_daemonxxLAST : std_logic_vector(0 downto 0);
    signal xxe_block_daemonxxNOT_LAST : std_logic_vector(0 downto 0);
    signal xxe_block_daemonxxRConstant_1 : std_logic_vector(7 downto 0);
    signal xxe_block_daemonxxZERO_COUNT : std_logic_vector(14 downto 0);
    -- 
  begin -- 
    R_LAST_13923_wire_constant <= "1";
    R_NOT_LAST_13851_wire_constant <= "0";
    R_NOT_LAST_13859_wire_constant <= "0";
    R_NOT_LAST_13867_wire_constant <= "0";
    R_NOT_LAST_13875_wire_constant <= "0";
    R_NOT_LAST_13883_wire_constant <= "0";
    R_NOT_LAST_13891_wire_constant <= "0";
    R_NOT_LAST_13899_wire_constant <= "0";
    R_NOT_LAST_13907_wire_constant <= "0";
    R_NOT_LAST_13915_wire_constant <= "0";
    R_RConstant_1_13773_wire_constant <= "00000001";
    R_ZERO_COUNT_13832_wire_constant <= "000000000000000";
    konst_13738_wire_constant <= "1";
    konst_13758_wire_constant <= "0";
    konst_13931_wire_constant <= "000000000000001";
    konst_13939_wire_constant <= "1";
    konst_13958_wire_constant <= "1";
    xxe_block_daemonxxLAST <= "1";
    xxe_block_daemonxxNOT_LAST <= "0";
    xxe_block_daemonxxRConstant_1 <= "00000001";
    xxe_block_daemonxxZERO_COUNT <= "000000000000000";
    phi_stmt_13763: Block -- phi operator 
      signal idata: std_logic_vector(255 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= e_init_key_13755_13765_buffered & e_new_key_13955_13766_buffered;
      req <= phi_stmt_13763_req_0 & phi_stmt_13763_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_13763",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 128) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_13763_ack_0,
          idata => idata,
          odata => K0_13763,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_13763
    phi_stmt_13767: Block -- phi operator 
      signal idata: std_logic_vector(29 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= e_init_count_13751_13769_buffered & e_new_count_13951_13770_buffered;
      req <= phi_stmt_13767_req_0 & phi_stmt_13767_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_13767",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 15) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_13767_ack_0,
          idata => idata,
          odata => countA_13767,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_13767
    phi_stmt_13823: Block -- phi operator 
      signal idata: std_logic_vector(29 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= countA_13767_13825_buffered & e_new_count_13951_13826_buffered;
      req <= phi_stmt_13823_req_0 & phi_stmt_13823_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_13823",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 15) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_13823_ack_0,
          idata => idata,
          odata => countB_13823,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_13823
    phi_stmt_13830: Block -- phi operator 
      signal idata: std_logic_vector(29 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_COUNT_13832_wire_constant & n_count_var_13933_13833_buffered;
      req <= phi_stmt_13830_req_0 & phi_stmt_13830_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_13830",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 15) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_13830_ack_0,
          idata => idata,
          odata => count_var_13830,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_13830
    -- flow-through slice operator slice_13746_inst
    e_get_key_13747 <= e_init_cmd_13743(143 downto 143);
    -- flow-through slice operator slice_13750_inst
    e_init_count_13751 <= e_init_cmd_13743(142 downto 128);
    -- flow-through slice operator slice_13754_inst
    e_init_key_13755 <= e_init_cmd_13743(127 downto 0);
    -- flow-through slice operator slice_13946_inst
    e_get_new_key_13947 <= e_new_cmd_13943(143 downto 143);
    -- flow-through slice operator slice_13950_inst
    e_new_count_13951 <= e_new_cmd_13943(142 downto 128);
    -- flow-through slice operator slice_13954_inst
    e_new_key_13955 <= e_new_cmd_13943(127 downto 0);
    W_K10_13856_delayed_10_13918_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_K10_13856_delayed_10_13918_inst_req_0;
      W_K10_13856_delayed_10_13918_inst_ack_0<= wack(0);
      rreq(0) <= W_K10_13856_delayed_10_13918_inst_req_1;
      W_K10_13856_delayed_10_13918_inst_ack_1<= rack(0);
      W_K10_13856_delayed_10_13918_inst : InterlockBuffer generic map ( -- 
        name => "W_K10_13856_delayed_10_13918_inst",
        buffer_size => 10,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 128,
        out_data_width => 128,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => K10_13821,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => K10_13856_delayed_10_13920,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_K1_13811_delayed_1_13846_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_K1_13811_delayed_1_13846_inst_req_0;
      W_K1_13811_delayed_1_13846_inst_ack_0<= wack(0);
      rreq(0) <= W_K1_13811_delayed_1_13846_inst_req_1;
      W_K1_13811_delayed_1_13846_inst_ack_1<= rack(0);
      W_K1_13811_delayed_1_13846_inst : InterlockBuffer generic map ( -- 
        name => "W_K1_13811_delayed_1_13846_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 128,
        out_data_width => 128,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => K1_13776,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => K1_13811_delayed_1_13848,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_K2_13816_delayed_2_13854_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_K2_13816_delayed_2_13854_inst_req_0;
      W_K2_13816_delayed_2_13854_inst_ack_0<= wack(0);
      rreq(0) <= W_K2_13816_delayed_2_13854_inst_req_1;
      W_K2_13816_delayed_2_13854_inst_ack_1<= rack(0);
      W_K2_13816_delayed_2_13854_inst : InterlockBuffer generic map ( -- 
        name => "W_K2_13816_delayed_2_13854_inst",
        buffer_size => 2,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 128,
        out_data_width => 128,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => K2_13781,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => K2_13816_delayed_2_13856,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_K3_13821_delayed_3_13862_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_K3_13821_delayed_3_13862_inst_req_0;
      W_K3_13821_delayed_3_13862_inst_ack_0<= wack(0);
      rreq(0) <= W_K3_13821_delayed_3_13862_inst_req_1;
      W_K3_13821_delayed_3_13862_inst_ack_1<= rack(0);
      W_K3_13821_delayed_3_13862_inst : InterlockBuffer generic map ( -- 
        name => "W_K3_13821_delayed_3_13862_inst",
        buffer_size => 3,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 128,
        out_data_width => 128,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => K3_13786,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => K3_13821_delayed_3_13864,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_K4_13826_delayed_4_13870_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_K4_13826_delayed_4_13870_inst_req_0;
      W_K4_13826_delayed_4_13870_inst_ack_0<= wack(0);
      rreq(0) <= W_K4_13826_delayed_4_13870_inst_req_1;
      W_K4_13826_delayed_4_13870_inst_ack_1<= rack(0);
      W_K4_13826_delayed_4_13870_inst : InterlockBuffer generic map ( -- 
        name => "W_K4_13826_delayed_4_13870_inst",
        buffer_size => 4,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 128,
        out_data_width => 128,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => K4_13791,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => K4_13826_delayed_4_13872,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_K5_13831_delayed_5_13878_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_K5_13831_delayed_5_13878_inst_req_0;
      W_K5_13831_delayed_5_13878_inst_ack_0<= wack(0);
      rreq(0) <= W_K5_13831_delayed_5_13878_inst_req_1;
      W_K5_13831_delayed_5_13878_inst_ack_1<= rack(0);
      W_K5_13831_delayed_5_13878_inst : InterlockBuffer generic map ( -- 
        name => "W_K5_13831_delayed_5_13878_inst",
        buffer_size => 5,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 128,
        out_data_width => 128,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => K5_13796,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => K5_13831_delayed_5_13880,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_K6_13836_delayed_6_13886_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_K6_13836_delayed_6_13886_inst_req_0;
      W_K6_13836_delayed_6_13886_inst_ack_0<= wack(0);
      rreq(0) <= W_K6_13836_delayed_6_13886_inst_req_1;
      W_K6_13836_delayed_6_13886_inst_ack_1<= rack(0);
      W_K6_13836_delayed_6_13886_inst : InterlockBuffer generic map ( -- 
        name => "W_K6_13836_delayed_6_13886_inst",
        buffer_size => 6,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 128,
        out_data_width => 128,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => K6_13801,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => K6_13836_delayed_6_13888,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_K7_13841_delayed_7_13894_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_K7_13841_delayed_7_13894_inst_req_0;
      W_K7_13841_delayed_7_13894_inst_ack_0<= wack(0);
      rreq(0) <= W_K7_13841_delayed_7_13894_inst_req_1;
      W_K7_13841_delayed_7_13894_inst_ack_1<= rack(0);
      W_K7_13841_delayed_7_13894_inst : InterlockBuffer generic map ( -- 
        name => "W_K7_13841_delayed_7_13894_inst",
        buffer_size => 7,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 128,
        out_data_width => 128,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => K7_13806,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => K7_13841_delayed_7_13896,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_K8_13846_delayed_8_13902_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_K8_13846_delayed_8_13902_inst_req_0;
      W_K8_13846_delayed_8_13902_inst_ack_0<= wack(0);
      rreq(0) <= W_K8_13846_delayed_8_13902_inst_req_1;
      W_K8_13846_delayed_8_13902_inst_ack_1<= rack(0);
      W_K8_13846_delayed_8_13902_inst : InterlockBuffer generic map ( -- 
        name => "W_K8_13846_delayed_8_13902_inst",
        buffer_size => 8,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 128,
        out_data_width => 128,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => K8_13811,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => K8_13846_delayed_8_13904,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_K9_13851_delayed_9_13910_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_K9_13851_delayed_9_13910_inst_req_0;
      W_K9_13851_delayed_9_13910_inst_ack_0<= wack(0);
      rreq(0) <= W_K9_13851_delayed_9_13910_inst_req_1;
      W_K9_13851_delayed_9_13910_inst_ack_1<= rack(0);
      W_K9_13851_delayed_9_13910_inst : InterlockBuffer generic map ( -- 
        name => "W_K9_13851_delayed_9_13910_inst",
        buffer_size => 9,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 128,
        out_data_width => 128,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => K9_13816,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => K9_13851_delayed_9_13912,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_round_S0_13810_delayed_1_13843_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_round_S0_13810_delayed_1_13843_inst_req_0;
      W_round_S0_13810_delayed_1_13843_inst_ack_0<= wack(0);
      rreq(0) <= W_round_S0_13810_delayed_1_13843_inst_req_1;
      W_round_S0_13810_delayed_1_13843_inst_ack_1<= rack(0);
      W_round_S0_13810_delayed_1_13843_inst : InterlockBuffer generic map ( -- 
        name => "W_round_S0_13810_delayed_1_13843_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 128,
        out_data_width => 128,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => round_S0_13842,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => round_S0_13810_delayed_1_13845,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    countA_13767_13825_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= countA_13767_13825_buf_req_0;
      countA_13767_13825_buf_ack_0<= wack(0);
      rreq(0) <= countA_13767_13825_buf_req_1;
      countA_13767_13825_buf_ack_1<= rack(0);
      countA_13767_13825_buf : InterlockBuffer generic map ( -- 
        name => "countA_13767_13825_buf",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 15,
        out_data_width => 15,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => countA_13767,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => countA_13767_13825_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    e_init_count_13751_13769_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= e_init_count_13751_13769_buf_req_0;
      e_init_count_13751_13769_buf_ack_0<= wack(0);
      rreq(0) <= e_init_count_13751_13769_buf_req_1;
      e_init_count_13751_13769_buf_ack_1<= rack(0);
      e_init_count_13751_13769_buf : InterlockBuffer generic map ( -- 
        name => "e_init_count_13751_13769_buf",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 15,
        out_data_width => 15,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => e_init_count_13751,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => e_init_count_13751_13769_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    e_init_key_13755_13765_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= e_init_key_13755_13765_buf_req_0;
      e_init_key_13755_13765_buf_ack_0<= wack(0);
      rreq(0) <= e_init_key_13755_13765_buf_req_1;
      e_init_key_13755_13765_buf_ack_1<= rack(0);
      e_init_key_13755_13765_buf : InterlockBuffer generic map ( -- 
        name => "e_init_key_13755_13765_buf",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 128,
        out_data_width => 128,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => e_init_key_13755,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => e_init_key_13755_13765_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    e_new_count_13951_13770_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= e_new_count_13951_13770_buf_req_0;
      e_new_count_13951_13770_buf_ack_0<= wack(0);
      rreq(0) <= e_new_count_13951_13770_buf_req_1;
      e_new_count_13951_13770_buf_ack_1<= rack(0);
      e_new_count_13951_13770_buf : InterlockBuffer generic map ( -- 
        name => "e_new_count_13951_13770_buf",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 15,
        out_data_width => 15,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => e_new_count_13951,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => e_new_count_13951_13770_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    e_new_count_13951_13826_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= e_new_count_13951_13826_buf_req_0;
      e_new_count_13951_13826_buf_ack_0<= wack(0);
      rreq(0) <= e_new_count_13951_13826_buf_req_1;
      e_new_count_13951_13826_buf_ack_1<= rack(0);
      e_new_count_13951_13826_buf : InterlockBuffer generic map ( -- 
        name => "e_new_count_13951_13826_buf",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 15,
        out_data_width => 15,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => e_new_count_13951,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => e_new_count_13951_13826_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    e_new_key_13955_13766_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= e_new_key_13955_13766_buf_req_0;
      e_new_key_13955_13766_buf_ack_0<= wack(0);
      rreq(0) <= e_new_key_13955_13766_buf_req_1;
      e_new_key_13955_13766_buf_ack_1<= rack(0);
      e_new_key_13955_13766_buf : InterlockBuffer generic map ( -- 
        name => "e_new_key_13955_13766_buf",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 128,
        out_data_width => 128,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => e_new_key_13955,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => e_new_key_13955_13766_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_count_var_13933_13833_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_count_var_13933_13833_buf_req_0;
      n_count_var_13933_13833_buf_ack_0<= wack(0);
      rreq(0) <= n_count_var_13933_13833_buf_req_1;
      n_count_var_13933_13833_buf_ack_1<= rack(0);
      n_count_var_13933_13833_buf : InterlockBuffer generic map ( -- 
        name => "n_count_var_13933_13833_buf",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 15,
        out_data_width => 15,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_count_var_13933,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_count_var_13933_13833_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    do_while_stmt_13828_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= ULT_u15_u1_13937_wire;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_13828_branch", condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_13828_branch_req_0,
          ack0 => do_while_stmt_13828_branch_ack_0,
          ack1 => do_while_stmt_13828_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_13756_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= EQ_u1_u1_13759_wire;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_13756_branch", condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_13756_branch_req_0,
          ack0 => if_stmt_13756_branch_ack_0,
          ack1 => if_stmt_13756_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_13956_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= EQ_u1_u1_13959_wire;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_13956_branch", condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_13956_branch_req_0,
          ack0 => if_stmt_13956_branch_ack_0,
          ack1 => if_stmt_13956_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- shared split operator group (0) : ADD_u15_u15_13932_inst 
    ApIntAdd_group_0: Block -- 
      signal data_in: std_logic_vector(14 downto 0);
      signal data_out: std_logic_vector(14 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= count_var_13830;
      n_count_var_13933 <= data_out(14 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u15_u15_13932_inst_req_0;
      ADD_u15_u15_13932_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u15_u15_13932_inst_req_1;
      ADD_u15_u15_13932_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(name => "gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_0",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 15,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 15,
          constant_operand => "000000000000001",
          constant_width => 15,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- binary operator EQ_u1_u1_13759_inst
    process(e_get_key_13747) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(e_get_key_13747, konst_13758_wire_constant, tmp_var);
      EQ_u1_u1_13759_wire <= tmp_var; -- 
    end process;
    -- binary operator EQ_u1_u1_13959_inst
    process(e_get_new_key_13947) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(e_get_new_key_13947, konst_13958_wire_constant, tmp_var);
      EQ_u1_u1_13959_wire <= tmp_var; -- 
    end process;
    -- binary operator ULT_u15_u1_13937_inst
    process(n_count_var_13933, countB_13823) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(n_count_var_13933, countB_13823, tmp_var);
      ULT_u15_u1_13937_wire <= tmp_var; -- 
    end process;
    -- binary operator XOR_u128_u128_13841_inst
    process(in128_13837, K0_13763) -- 
      variable tmp_var : std_logic_vector(127 downto 0); -- 
    begin -- 
      ApIntXor_proc(in128_13837, K0_13763, tmp_var);
      round_S0_13842 <= tmp_var; -- 
    end process;
    -- shared inport operator group (0) : RPIPE_e_cmd_pipe_13742_inst RPIPE_e_cmd_pipe_13942_inst 
    InportGroup0: Block -- 
      signal data_out: std_logic_vector(287 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 1 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= RPIPE_e_cmd_pipe_13742_inst_req_0;
      reqL_unguarded(0) <= RPIPE_e_cmd_pipe_13942_inst_req_0;
      RPIPE_e_cmd_pipe_13742_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_e_cmd_pipe_13942_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= RPIPE_e_cmd_pipe_13742_inst_req_1;
      reqR_unguarded(0) <= RPIPE_e_cmd_pipe_13942_inst_req_1;
      RPIPE_e_cmd_pipe_13742_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_e_cmd_pipe_13942_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      gI: SplitGuardInterface generic map(name => "gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      e_init_cmd_13743 <= data_out(287 downto 144);
      e_new_cmd_13943 <= data_out(143 downto 0);
      e_cmd_pipe_read_0: InputPortRevised -- 
        generic map ( name => "e_cmd_pipe_read_0", data_width => 144,  num_reqs => 2,  output_buffering => outBUFs,   no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => e_cmd_pipe_pipe_read_req(0),
          oack => e_cmd_pipe_pipe_read_ack(0),
          odata => e_cmd_pipe_pipe_read_data(143 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared inport operator group (1) : RPIPE_e_in_buf_13836_inst 
    InportGroup1: Block -- 
      signal data_out: std_logic_vector(127 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_e_in_buf_13836_inst_req_0;
      RPIPE_e_in_buf_13836_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_e_in_buf_13836_inst_req_1;
      RPIPE_e_in_buf_13836_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      gI: SplitGuardInterface generic map(name => "gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      in128_13837 <= data_out(127 downto 0);
      e_in_buf_read_1: InputPortRevised -- 
        generic map ( name => "e_in_buf_read_1", data_width => 128,  num_reqs => 1,  output_buffering => outBUFs,   no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => e_in_buf_pipe_read_req(0),
          oack => e_in_buf_pipe_read_ack(0),
          odata => e_in_buf_pipe_read_data(127 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 1
    -- shared outport operator group (0) : WPIPE_e_block_done_13737_inst WPIPE_e_block_done_13938_inst 
    OutportGroup0: Block -- 
      signal data_in: std_logic_vector(1 downto 0);
      signal sample_req, sample_ack : BooleanArray( 1 downto 0);
      signal update_req, update_ack : BooleanArray( 1 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 1 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      sample_req_unguarded(1) <= WPIPE_e_block_done_13737_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_e_block_done_13938_inst_req_0;
      WPIPE_e_block_done_13737_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_e_block_done_13938_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(1) <= WPIPE_e_block_done_13737_inst_req_1;
      update_req_unguarded(0) <= WPIPE_e_block_done_13938_inst_req_1;
      WPIPE_e_block_done_13737_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_e_block_done_13938_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      gI: SplitGuardInterface generic map(name => "gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      data_in <= konst_13738_wire_constant & konst_13939_wire_constant;
      e_block_done_write_0: OutputPortRevised -- 
        generic map ( name => "e_block_done", data_width => 1, num_reqs => 2, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => e_block_done_pipe_write_req(0),
          oack => e_block_done_pipe_write_ack(0),
          odata => e_block_done_pipe_write_data(0 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_e_out_buf_13926_inst 
    OutportGroup1: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_e_out_buf_13926_inst_req_0;
      WPIPE_e_out_buf_13926_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_e_out_buf_13926_inst_req_1;
      WPIPE_e_out_buf_13926_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      gI: SplitGuardInterface generic map(name => "gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      data_in <= round_S10_13925;
      e_out_buf_write_1: OutputPortRevised -- 
        generic map ( name => "e_out_buf", data_width => 128, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => e_out_buf_pipe_write_req(0),
          oack => e_out_buf_pipe_write_ack(0),
          odata => e_out_buf_pipe_write_data(127 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared call operator group (0) : call_stmt_13781_call call_stmt_13776_call call_stmt_13821_call call_stmt_13816_call call_stmt_13811_call call_stmt_13806_call call_stmt_13801_call call_stmt_13796_call call_stmt_13791_call call_stmt_13786_call 
    key_expand_single_call_group_0: Block -- 
      signal data_in: std_logic_vector(1359 downto 0);
      signal data_out: std_logic_vector(1359 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 9 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 9 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 9 downto 0);
      signal guard_vector : std_logic_vector( 9 downto 0);
      constant inBUFs : IntegerArray(9 downto 0) := (9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(9 downto 0) := (9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(9 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false);
      constant guardBuffering: IntegerArray(9 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2);
      -- 
    begin -- 
      reqL_unguarded(9) <= call_stmt_13781_call_req_0;
      reqL_unguarded(8) <= call_stmt_13776_call_req_0;
      reqL_unguarded(7) <= call_stmt_13821_call_req_0;
      reqL_unguarded(6) <= call_stmt_13816_call_req_0;
      reqL_unguarded(5) <= call_stmt_13811_call_req_0;
      reqL_unguarded(4) <= call_stmt_13806_call_req_0;
      reqL_unguarded(3) <= call_stmt_13801_call_req_0;
      reqL_unguarded(2) <= call_stmt_13796_call_req_0;
      reqL_unguarded(1) <= call_stmt_13791_call_req_0;
      reqL_unguarded(0) <= call_stmt_13786_call_req_0;
      call_stmt_13781_call_ack_0 <= ackL_unguarded(9);
      call_stmt_13776_call_ack_0 <= ackL_unguarded(8);
      call_stmt_13821_call_ack_0 <= ackL_unguarded(7);
      call_stmt_13816_call_ack_0 <= ackL_unguarded(6);
      call_stmt_13811_call_ack_0 <= ackL_unguarded(5);
      call_stmt_13806_call_ack_0 <= ackL_unguarded(4);
      call_stmt_13801_call_ack_0 <= ackL_unguarded(3);
      call_stmt_13796_call_ack_0 <= ackL_unguarded(2);
      call_stmt_13791_call_ack_0 <= ackL_unguarded(1);
      call_stmt_13786_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(9) <= call_stmt_13781_call_req_1;
      reqR_unguarded(8) <= call_stmt_13776_call_req_1;
      reqR_unguarded(7) <= call_stmt_13821_call_req_1;
      reqR_unguarded(6) <= call_stmt_13816_call_req_1;
      reqR_unguarded(5) <= call_stmt_13811_call_req_1;
      reqR_unguarded(4) <= call_stmt_13806_call_req_1;
      reqR_unguarded(3) <= call_stmt_13801_call_req_1;
      reqR_unguarded(2) <= call_stmt_13796_call_req_1;
      reqR_unguarded(1) <= call_stmt_13791_call_req_1;
      reqR_unguarded(0) <= call_stmt_13786_call_req_1;
      call_stmt_13781_call_ack_1 <= ackR_unguarded(9);
      call_stmt_13776_call_ack_1 <= ackR_unguarded(8);
      call_stmt_13821_call_ack_1 <= ackR_unguarded(7);
      call_stmt_13816_call_ack_1 <= ackR_unguarded(6);
      call_stmt_13811_call_ack_1 <= ackR_unguarded(5);
      call_stmt_13806_call_ack_1 <= ackR_unguarded(4);
      call_stmt_13801_call_ack_1 <= ackR_unguarded(3);
      call_stmt_13796_call_ack_1 <= ackR_unguarded(2);
      call_stmt_13791_call_ack_1 <= ackR_unguarded(1);
      call_stmt_13786_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      key_expand_single_call_group_0_accessRegulator_0: access_regulator_base generic map (name => "key_expand_single_call_group_0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      key_expand_single_call_group_0_accessRegulator_1: access_regulator_base generic map (name => "key_expand_single_call_group_0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      key_expand_single_call_group_0_accessRegulator_2: access_regulator_base generic map (name => "key_expand_single_call_group_0_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      key_expand_single_call_group_0_accessRegulator_3: access_regulator_base generic map (name => "key_expand_single_call_group_0_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      key_expand_single_call_group_0_accessRegulator_4: access_regulator_base generic map (name => "key_expand_single_call_group_0_accessRegulator_4", num_slots => 1) -- 
        port map (req => reqL_unregulated(4), -- 
          ack => ackL_unregulated(4),
          regulated_req => reqL(4),
          regulated_ack => ackL(4),
          release_req => reqR(4),
          release_ack => ackR(4),
          clk => clk, reset => reset); -- 
      key_expand_single_call_group_0_accessRegulator_5: access_regulator_base generic map (name => "key_expand_single_call_group_0_accessRegulator_5", num_slots => 1) -- 
        port map (req => reqL_unregulated(5), -- 
          ack => ackL_unregulated(5),
          regulated_req => reqL(5),
          regulated_ack => ackL(5),
          release_req => reqR(5),
          release_ack => ackR(5),
          clk => clk, reset => reset); -- 
      key_expand_single_call_group_0_accessRegulator_6: access_regulator_base generic map (name => "key_expand_single_call_group_0_accessRegulator_6", num_slots => 1) -- 
        port map (req => reqL_unregulated(6), -- 
          ack => ackL_unregulated(6),
          regulated_req => reqL(6),
          regulated_ack => ackL(6),
          release_req => reqR(6),
          release_ack => ackR(6),
          clk => clk, reset => reset); -- 
      key_expand_single_call_group_0_accessRegulator_7: access_regulator_base generic map (name => "key_expand_single_call_group_0_accessRegulator_7", num_slots => 1) -- 
        port map (req => reqL_unregulated(7), -- 
          ack => ackL_unregulated(7),
          regulated_req => reqL(7),
          regulated_ack => ackL(7),
          release_req => reqR(7),
          release_ack => ackR(7),
          clk => clk, reset => reset); -- 
      key_expand_single_call_group_0_accessRegulator_8: access_regulator_base generic map (name => "key_expand_single_call_group_0_accessRegulator_8", num_slots => 1) -- 
        port map (req => reqL_unregulated(8), -- 
          ack => ackL_unregulated(8),
          regulated_req => reqL(8),
          regulated_ack => ackL(8),
          release_req => reqR(8),
          release_ack => ackR(8),
          clk => clk, reset => reset); -- 
      key_expand_single_call_group_0_accessRegulator_9: access_regulator_base generic map (name => "key_expand_single_call_group_0_accessRegulator_9", num_slots => 1) -- 
        port map (req => reqL_unregulated(9), -- 
          ack => ackL_unregulated(9),
          regulated_req => reqL(9),
          regulated_ack => ackL(9),
          release_req => reqR(9),
          release_ack => ackR(9),
          clk => clk, reset => reset); -- 
      gI: SplitGuardInterface generic map(name => "gI", nreqs => 10, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= K1_13776 & RConstant_2_13776 & K0_13763 & R_RConstant_1_13773_wire_constant & K9_13816 & RConstant_10_13816 & K8_13811 & RConstant_9_13811 & K7_13806 & RConstant_8_13806 & K6_13801 & RConstant_7_13801 & K5_13796 & RConstant_6_13796 & K4_13791 & RConstant_5_13791 & K3_13786 & RConstant_4_13786 & K2_13781 & RConstant_3_13781;
      K2_13781 <= data_out(1359 downto 1232);
      RConstant_3_13781 <= data_out(1231 downto 1224);
      K1_13776 <= data_out(1223 downto 1096);
      RConstant_2_13776 <= data_out(1095 downto 1088);
      K10_13821 <= data_out(1087 downto 960);
      RConstant_11_13821 <= data_out(959 downto 952);
      K9_13816 <= data_out(951 downto 824);
      RConstant_10_13816 <= data_out(823 downto 816);
      K8_13811 <= data_out(815 downto 688);
      RConstant_9_13811 <= data_out(687 downto 680);
      K7_13806 <= data_out(679 downto 552);
      RConstant_8_13806 <= data_out(551 downto 544);
      K6_13801 <= data_out(543 downto 416);
      RConstant_7_13801 <= data_out(415 downto 408);
      K5_13796 <= data_out(407 downto 280);
      RConstant_6_13796 <= data_out(279 downto 272);
      K4_13791 <= data_out(271 downto 144);
      RConstant_5_13791 <= data_out(143 downto 136);
      K3_13786 <= data_out(135 downto 8);
      RConstant_4_13786 <= data_out(7 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 1360,
        owidth => 136,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 4,
        nreqs => 10,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => key_expand_single_call_reqs(0),
          ackR => key_expand_single_call_acks(0),
          dataR => key_expand_single_call_data(135 downto 0),
          tagR => key_expand_single_call_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 136,
          owidth => 1360,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 4,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 10) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => key_expand_single_return_acks(0), -- cross-over
          ackL => key_expand_single_return_reqs(0), -- cross-over
          dataL => key_expand_single_return_data(135 downto 0),
          tagL => key_expand_single_return_tag(3 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    call_stmt_13853_call_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= call_stmt_13853_call_req_0;
      call_stmt_13853_call_ack_0<= sample_ack(0);
      update_req(0) <= call_stmt_13853_call_req_1;
      call_stmt_13853_call_ack_1<= update_ack(0);
      call_stmt_13853_call: enc_round_Operator  port map ( -- 
        sample_req => sample_req(0), 
        sample_ack => sample_ack(0), 
        update_req => update_req(0), 
        update_ack => update_ack(0), 
        round_in => round_S0_13810_delayed_1_13845,
        key_in => K1_13811_delayed_1_13848,
        l_round => R_NOT_LAST_13851_wire_constant,
        round_out => round_S1_13853,
        clk => clk, reset => reset  
        -- 
      );-- 
    end block;
    call_stmt_13861_call_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= call_stmt_13861_call_req_0;
      call_stmt_13861_call_ack_0<= sample_ack(0);
      update_req(0) <= call_stmt_13861_call_req_1;
      call_stmt_13861_call_ack_1<= update_ack(0);
      call_stmt_13861_call: enc_round_Operator  port map ( -- 
        sample_req => sample_req(0), 
        sample_ack => sample_ack(0), 
        update_req => update_req(0), 
        update_ack => update_ack(0), 
        round_in => round_S1_13853,
        key_in => K2_13816_delayed_2_13856,
        l_round => R_NOT_LAST_13859_wire_constant,
        round_out => round_S2_13861,
        clk => clk, reset => reset  
        -- 
      );-- 
    end block;
    call_stmt_13869_call_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= call_stmt_13869_call_req_0;
      call_stmt_13869_call_ack_0<= sample_ack(0);
      update_req(0) <= call_stmt_13869_call_req_1;
      call_stmt_13869_call_ack_1<= update_ack(0);
      call_stmt_13869_call: enc_round_Operator  port map ( -- 
        sample_req => sample_req(0), 
        sample_ack => sample_ack(0), 
        update_req => update_req(0), 
        update_ack => update_ack(0), 
        round_in => round_S2_13861,
        key_in => K3_13821_delayed_3_13864,
        l_round => R_NOT_LAST_13867_wire_constant,
        round_out => round_S3_13869,
        clk => clk, reset => reset  
        -- 
      );-- 
    end block;
    call_stmt_13877_call_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= call_stmt_13877_call_req_0;
      call_stmt_13877_call_ack_0<= sample_ack(0);
      update_req(0) <= call_stmt_13877_call_req_1;
      call_stmt_13877_call_ack_1<= update_ack(0);
      call_stmt_13877_call: enc_round_Operator  port map ( -- 
        sample_req => sample_req(0), 
        sample_ack => sample_ack(0), 
        update_req => update_req(0), 
        update_ack => update_ack(0), 
        round_in => round_S3_13869,
        key_in => K4_13826_delayed_4_13872,
        l_round => R_NOT_LAST_13875_wire_constant,
        round_out => round_S4_13877,
        clk => clk, reset => reset  
        -- 
      );-- 
    end block;
    call_stmt_13885_call_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= call_stmt_13885_call_req_0;
      call_stmt_13885_call_ack_0<= sample_ack(0);
      update_req(0) <= call_stmt_13885_call_req_1;
      call_stmt_13885_call_ack_1<= update_ack(0);
      call_stmt_13885_call: enc_round_Operator  port map ( -- 
        sample_req => sample_req(0), 
        sample_ack => sample_ack(0), 
        update_req => update_req(0), 
        update_ack => update_ack(0), 
        round_in => round_S4_13877,
        key_in => K5_13831_delayed_5_13880,
        l_round => R_NOT_LAST_13883_wire_constant,
        round_out => round_S5_13885,
        clk => clk, reset => reset  
        -- 
      );-- 
    end block;
    call_stmt_13893_call_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= call_stmt_13893_call_req_0;
      call_stmt_13893_call_ack_0<= sample_ack(0);
      update_req(0) <= call_stmt_13893_call_req_1;
      call_stmt_13893_call_ack_1<= update_ack(0);
      call_stmt_13893_call: enc_round_Operator  port map ( -- 
        sample_req => sample_req(0), 
        sample_ack => sample_ack(0), 
        update_req => update_req(0), 
        update_ack => update_ack(0), 
        round_in => round_S5_13885,
        key_in => K6_13836_delayed_6_13888,
        l_round => R_NOT_LAST_13891_wire_constant,
        round_out => round_S6_13893,
        clk => clk, reset => reset  
        -- 
      );-- 
    end block;
    call_stmt_13901_call_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= call_stmt_13901_call_req_0;
      call_stmt_13901_call_ack_0<= sample_ack(0);
      update_req(0) <= call_stmt_13901_call_req_1;
      call_stmt_13901_call_ack_1<= update_ack(0);
      call_stmt_13901_call: enc_round_Operator  port map ( -- 
        sample_req => sample_req(0), 
        sample_ack => sample_ack(0), 
        update_req => update_req(0), 
        update_ack => update_ack(0), 
        round_in => round_S6_13893,
        key_in => K7_13841_delayed_7_13896,
        l_round => R_NOT_LAST_13899_wire_constant,
        round_out => round_S7_13901,
        clk => clk, reset => reset  
        -- 
      );-- 
    end block;
    call_stmt_13909_call_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= call_stmt_13909_call_req_0;
      call_stmt_13909_call_ack_0<= sample_ack(0);
      update_req(0) <= call_stmt_13909_call_req_1;
      call_stmt_13909_call_ack_1<= update_ack(0);
      call_stmt_13909_call: enc_round_Operator  port map ( -- 
        sample_req => sample_req(0), 
        sample_ack => sample_ack(0), 
        update_req => update_req(0), 
        update_ack => update_ack(0), 
        round_in => round_S7_13901,
        key_in => K8_13846_delayed_8_13904,
        l_round => R_NOT_LAST_13907_wire_constant,
        round_out => round_S8_13909,
        clk => clk, reset => reset  
        -- 
      );-- 
    end block;
    call_stmt_13917_call_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= call_stmt_13917_call_req_0;
      call_stmt_13917_call_ack_0<= sample_ack(0);
      update_req(0) <= call_stmt_13917_call_req_1;
      call_stmt_13917_call_ack_1<= update_ack(0);
      call_stmt_13917_call: enc_round_Operator  port map ( -- 
        sample_req => sample_req(0), 
        sample_ack => sample_ack(0), 
        update_req => update_req(0), 
        update_ack => update_ack(0), 
        round_in => round_S8_13909,
        key_in => K9_13851_delayed_9_13912,
        l_round => R_NOT_LAST_13915_wire_constant,
        round_out => round_S9_13917,
        clk => clk, reset => reset  
        -- 
      );-- 
    end block;
    call_stmt_13925_call_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= call_stmt_13925_call_req_0;
      call_stmt_13925_call_ack_0<= sample_ack(0);
      update_req(0) <= call_stmt_13925_call_req_1;
      call_stmt_13925_call_ack_1<= update_ack(0);
      call_stmt_13925_call: enc_round_Operator  port map ( -- 
        sample_req => sample_req(0), 
        sample_ack => sample_ack(0), 
        update_req => update_req(0), 
        update_ack => update_ack(0), 
        round_in => round_S9_13917,
        key_in => K10_13856_delayed_10_13920,
        l_round => R_LAST_13923_wire_constant,
        round_out => round_S10_13925,
        clk => clk, reset => reset  
        -- 
      );-- 
    end block;
    -- 
  end Block; -- data_path
  -- 
end e_block_daemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library work;
use work.ahir_system_global_package.all;
entity enc_round_Operator is -- 
  port ( -- 
    sample_req: in boolean;
    sample_ack: out boolean;
    update_req: in boolean;
    update_ack: out boolean;
    round_in : in  std_logic_vector(127 downto 0);
    key_in : in  std_logic_vector(127 downto 0);
    l_round : in  std_logic_vector(0 downto 0);
    round_out : out  std_logic_vector(127 downto 0);
    clk, reset: in std_logic
    -- 
  );
  -- 
end entity enc_round_Operator;
architecture enc_round_Operator_arch of enc_round_Operator is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal update_ack_symbol: Boolean;
  signal default_zero_sig: std_logic;
  -- input port buffer signals
  signal round_in_buffer :  std_logic_vector(127 downto 0);
  signal round_in_update_enable: Boolean;
  signal round_in_update_enable_unmarked: Boolean;
  signal key_in_buffer :  std_logic_vector(127 downto 0);
  signal key_in_update_enable: Boolean;
  signal key_in_update_enable_unmarked: Boolean;
  signal l_round_buffer :  std_logic_vector(0 downto 0);
  signal l_round_update_enable: Boolean;
  signal l_round_update_enable_unmarked: Boolean;
  -- output port buffer signals
  signal round_out_buffer :  std_logic_vector(127 downto 0);
  signal round_out_update_enable: Boolean;
  signal enc_round_CP_7671_start: Boolean;
  signal enc_round_CP_7671_symbol: Boolean;
  signal cp_all_inputs_sampled: Boolean;
  -- volatile/operator module components. 
  component sbox_mux_impl_Volatile is -- 
    port ( -- 
      data_in : in  std_logic_vector(7 downto 0);
      s_out : out  std_logic_vector(7 downto 0)-- 
    );
    -- 
  end component; 
  -- links between control-path and data-path
  signal XOR_u128_u128_13720_inst_req_0 : boolean;
  signal XOR_u128_u128_13720_inst_ack_0 : boolean;
  signal XOR_u128_u128_13720_inst_req_1 : boolean;
  signal XOR_u128_u128_13720_inst_ack_1 : boolean;
  -- 
begin --  
  sample_ack <= enc_round_CP_7671_symbol;
  -- input handling ------------------------------------------------
  round_in_buffer <= round_in;
  key_in_buffer <= key_in;
  l_round_buffer <= l_round;
  enc_round_CP_7671_start <= sample_req;
  -- output handling  -------------------------------------------------------
  round_out <= round_out_buffer;
  round_out_update_enable <= update_req;
  update_ack_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 22) := "update_ack_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= enc_round_CP_7671_symbol & update_req;
    gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => update_ack_symbol, clk => clk, reset => reset); --
  end block;
  -- update ack. 
  update_ack <= update_ack_symbol;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  enc_round_CP_7671: Block -- control-path 
    signal enc_round_CP_7671_elements: BooleanArray(2 downto 0);
    -- 
  begin -- 
    enc_round_CP_7671_elements(0) <= enc_round_CP_7671_start;
    enc_round_CP_7671_symbol <= enc_round_CP_7671_elements(2);
    -- CP-element group 0:  join  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (3072) 
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13099_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13099_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13099_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Sa_13094_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13099_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13095_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13099_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13095_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13095_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13095_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13095_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Sa_13094_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13095_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13099_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13099_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Sa_13094_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13095_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13091_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Sa_13094_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Sb_13110_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Sb_13110_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13095_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13095_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13095_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13095_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13099_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13095_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Sb_13118_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Sb_13118_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Sb_13118_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Sb_13118_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13103_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13103_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13115_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13115_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13115_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13111_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Sa_13102_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13103_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13099_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13107_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13107_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13111_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13111_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Sa_13102_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Sa_13102_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Sa_13098_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13099_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13103_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13103_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13111_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13103_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Sa_13102_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Sa_13098_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13099_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13103_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13103_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13111_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13111_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13111_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13103_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13103_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Sa_13098_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13099_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13103_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13103_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13119_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13119_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13119_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13119_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13115_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Sb_13114_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Sb_13114_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13115_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13115_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13115_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Sd_13138_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Sd_13138_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13299_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13139_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Sb_13114_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Sb_13114_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Sc_13122_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Sc_13122_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Sc_13122_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13123_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13119_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13119_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13119_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13119_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13111_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S03x2_13315_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13115_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13115_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13115_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13294_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13119_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13119_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13119_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13119_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S02x2_13305_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Sb_13110_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Sb_13110_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13135_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13135_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13135_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S03x2_13318_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13111_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13111_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13115_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13115_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13123_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13123_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13123_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13123_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Sc_13122_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13111_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13111_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13135_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13135_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13135_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13135_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13135_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13107_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13299_complete/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Sc_13134_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Sc_13134_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Sc_13134_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13299_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13299_start/ack
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13299_start/req
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S01_13292_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13107_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13107_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13107_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13135_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13135_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13135_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13135_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Sc_13134_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13107_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13131_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13131_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13131_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13131_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13131_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13131_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13107_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13107_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13131_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Sc_13130_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Sc_13130_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Sc_13130_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Sc_13130_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S02_13302_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13131_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13131_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13107_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13127_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13127_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13127_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13127_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S03x2_13315_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13131_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13131_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13131_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Sb_13106_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Sb_13106_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Sc_13126_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Sc_13126_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Sc_13126_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S02_13302_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13127_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13127_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13127_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13127_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Sb_13106_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Sb_13106_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13123_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13123_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S03x2_13315_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13127_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13127_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13127_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13127_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Sc_13126_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13107_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13107_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13139_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13139_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13139_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13139_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Sd_13138_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Sd_13138_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13123_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13123_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13123_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13123_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13123_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/call_stmt_13176_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/call_stmt_13176_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13289_start/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13299_complete/req
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13307_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S00x2_13288_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S03x2_13318_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13307_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13289_start/req
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13304_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13329_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13329_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13314_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13304_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13294_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13294_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13294_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13299_complete/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13309_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13297_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13289_start/ack
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S02x2_13305_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S00x2_13288_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13299_complete/ack
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13299_start/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13289_complete/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13307_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13297_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13297_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13294_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13317_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13317_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S02x2_13305_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13319_start/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13289_complete/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S02_13302_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13294_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13289_start/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13319_start/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S01_13292_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13317_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13317_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13289_complete/req
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13289_complete/ack
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S00x2_13288_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S02x2_13305_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S01_13292_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S01_13292_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13319_start/req
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13319_start/ack
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S03x2_13318_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S03x2_13318_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13304_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13294_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13309_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13299_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13317_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13317_Update/$exit
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13299_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13297_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13075_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13075_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13075_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13075_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_round_in_13074_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_round_in_13074_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_round_in_13074_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_round_in_13074_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13075_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13075_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13075_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13075_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13075_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13075_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13075_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13075_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13079_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13079_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13079_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13079_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_round_in_13078_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_round_in_13078_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_round_in_13078_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_round_in_13078_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13079_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13079_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13079_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13079_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13079_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13079_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13079_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13079_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13083_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13083_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13083_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13083_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_round_in_13082_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_round_in_13082_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_round_in_13082_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_round_in_13082_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13083_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13083_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13083_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13083_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13083_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13083_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13083_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13083_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13087_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13087_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13087_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Sa_13098_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13087_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_round_in_13086_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_round_in_13086_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_round_in_13086_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_round_in_13086_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13087_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13087_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13087_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13087_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13087_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13087_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13087_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13087_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13091_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13091_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13091_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13091_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Sa_13090_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Sa_13090_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Sa_13090_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Sa_13090_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13091_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13091_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13091_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13091_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13091_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13091_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13091_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13139_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13139_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13139_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13139_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13139_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13139_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13139_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13143_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13143_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13143_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13143_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Sd_13142_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Sd_13142_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Sd_13142_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Sd_13142_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13143_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13143_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13143_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13143_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13143_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13143_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13143_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13143_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13147_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13147_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13147_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13147_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Sd_13146_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Sd_13146_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Sd_13146_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Sd_13146_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13147_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13147_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13147_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13147_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13147_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13147_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13147_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13147_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13151_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13151_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13151_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13151_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Sd_13150_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Sd_13150_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Sd_13150_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Sd_13150_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13151_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13151_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13151_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13151_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13151_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13151_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13151_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/slice_13151_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/call_stmt_13155_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/call_stmt_13155_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/call_stmt_13155_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/call_stmt_13155_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S00sr_13153_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S00sr_13153_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S00sr_13153_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S00sr_13153_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/call_stmt_13158_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/call_stmt_13158_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/call_stmt_13158_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/call_stmt_13158_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S05sr_13156_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S05sr_13156_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S05sr_13156_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S05sr_13156_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/call_stmt_13161_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/call_stmt_13161_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/call_stmt_13161_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/call_stmt_13161_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S10sr_13159_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S10sr_13159_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S10sr_13159_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S10sr_13159_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/call_stmt_13164_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/call_stmt_13164_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/call_stmt_13164_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/call_stmt_13164_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S15sr_13162_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S15sr_13162_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S15sr_13162_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S15sr_13162_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/call_stmt_13167_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/call_stmt_13167_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/call_stmt_13167_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/call_stmt_13167_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S04sr_13165_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S04sr_13165_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S04sr_13165_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S04sr_13165_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/call_stmt_13170_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/call_stmt_13170_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/call_stmt_13170_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/call_stmt_13170_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S09sr_13168_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S09sr_13168_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S09sr_13168_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S09sr_13168_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/call_stmt_13173_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/call_stmt_13173_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/call_stmt_13173_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/call_stmt_13173_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S14sr_13171_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S14sr_13171_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S14sr_13171_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S14sr_13171_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/call_stmt_13176_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13324_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13324_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13324_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13324_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S04_13322_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/call_stmt_13176_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S03sr_13174_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S03sr_13174_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S03sr_13174_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S03sr_13174_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/call_stmt_13179_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/call_stmt_13179_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/call_stmt_13179_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/call_stmt_13179_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S08sr_13177_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S08sr_13177_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S08sr_13177_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S08sr_13177_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/call_stmt_13182_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/call_stmt_13182_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/call_stmt_13182_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/call_stmt_13182_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S13sr_13180_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S13sr_13180_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S13sr_13180_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S13sr_13180_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/call_stmt_13185_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/call_stmt_13185_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/call_stmt_13185_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/call_stmt_13185_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S02sr_13183_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S02sr_13183_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S02sr_13183_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S02sr_13183_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/call_stmt_13188_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/call_stmt_13188_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/call_stmt_13188_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/call_stmt_13188_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S07sr_13186_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S07sr_13186_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S07sr_13186_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S07sr_13186_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/call_stmt_13191_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/call_stmt_13191_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/call_stmt_13191_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/call_stmt_13191_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S12sr_13189_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S12sr_13189_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S12sr_13189_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S12sr_13189_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S02_13302_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S03_13312_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S03_13312_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S03_13312_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/call_stmt_13194_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/call_stmt_13194_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/call_stmt_13194_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/call_stmt_13194_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13304_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S03x2_13315_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13317_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S01sr_13192_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S01sr_13192_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S01sr_13192_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S01sr_13192_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13304_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S03_13312_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13314_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13314_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13314_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/call_stmt_13197_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/call_stmt_13197_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/call_stmt_13197_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/call_stmt_13197_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13304_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13317_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13317_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S06sr_13195_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S06sr_13195_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S06sr_13195_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S06sr_13195_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13304_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13314_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13319_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13319_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13319_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/call_stmt_13200_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/call_stmt_13200_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/call_stmt_13200_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/call_stmt_13200_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13309_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13317_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13314_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S11sr_13198_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S11sr_13198_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S11sr_13198_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S11sr_13198_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13309_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13319_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13309_complete/ack
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13309_complete/req
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13309_complete/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13204_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13204_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13204_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13204_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S00_13202_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S00_13202_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S00_13202_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S00_13202_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13307_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13309_complete/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13309_start/ack
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13309_start/req
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13204_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13204_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13297_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13204_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13204_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13204_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13204_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13297_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13204_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13204_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13309_start/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13314_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13329_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13329_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13314_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13314_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13209_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13209_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13209_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13209_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S01_13207_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S01_13207_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S01_13207_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S01_13207_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13307_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13309_start/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S02x2_13308_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S02x2_13308_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13209_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13209_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13297_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13209_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13209_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13209_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13209_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S01x2_13295_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13209_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13209_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S02x2_13308_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13319_complete/req
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13319_complete/ack
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13314_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13314_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13214_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13214_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13214_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13214_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S02_13212_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S02_13212_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S02_13212_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S02_13212_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13307_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S02x2_13308_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13307_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13307_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13307_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13214_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13214_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S01x2_13295_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13214_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13214_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13214_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13214_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S01x2_13295_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13214_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13214_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13307_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13314_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13319_complete/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13319_complete/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13299_start/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13304_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13219_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13219_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13219_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13219_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S03_13217_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S03_13217_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S03_13217_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S03_13217_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13304_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13437_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13219_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13219_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S01x2_13295_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13219_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13219_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13219_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13219_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13297_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13219_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13219_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S01x2_13298_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S01x2_13298_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13304_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13224_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13224_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13224_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13224_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S04_13222_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S04_13222_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S04_13222_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S04_13222_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13304_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13448_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13437_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13224_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13224_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13297_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13224_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13224_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13224_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13224_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13297_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13224_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13224_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S01x2_13298_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13317_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S01x2_13298_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13229_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13229_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13229_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13229_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S05_13227_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S05_13227_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S05_13227_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S05_13227_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13304_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S15x2_13438_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13229_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13229_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13297_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13229_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13229_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13229_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13229_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13294_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13229_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13229_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13297_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13317_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13437_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13234_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13234_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13234_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13234_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S06_13232_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S06_13232_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S06_13232_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S06_13232_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13437_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13437_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13234_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13234_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13294_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13234_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13234_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13234_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13234_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13294_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13234_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13234_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13307_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13239_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13239_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13239_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13239_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S07_13237_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S07_13237_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S07_13237_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S07_13237_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13239_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13239_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13294_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13239_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13239_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13239_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13239_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13294_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13239_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13239_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13307_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13437_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13244_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13244_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13244_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13244_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S08_13242_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S08_13242_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S08_13242_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S08_13242_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S15x2_13438_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13437_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13244_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13244_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13244_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13244_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13244_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13244_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13244_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13244_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13457_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S15x2_13438_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13249_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13249_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13249_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13249_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S09_13247_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S09_13247_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S09_13247_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S09_13247_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13448_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13249_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13249_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13249_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13249_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13249_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13249_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13249_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13249_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13254_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13254_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13254_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13254_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S10_13252_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S10_13252_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S10_13252_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S10_13252_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13448_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S03_13446_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13448_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13254_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13254_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13254_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13254_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13254_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13254_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S00_13442_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13254_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13254_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S01_13443_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13259_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13259_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13259_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13259_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S11_13257_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S11_13257_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S11_13257_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S11_13257_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13448_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13457_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13259_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13259_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S00_13442_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13259_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13259_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13259_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13259_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S00_13442_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13259_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13259_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S15x2_13438_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S04_13451_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S04_13451_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13264_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13264_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13264_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13264_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S12_13262_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S12_13262_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S12_13262_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S12_13262_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13264_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13264_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13264_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13264_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13264_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13264_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S00_13442_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13264_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13264_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S03_13446_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S03_13446_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13453_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13437_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13269_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13269_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13269_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13269_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S13_13267_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S13_13267_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S13_13267_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S13_13267_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13448_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13269_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13269_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13269_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13269_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13269_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13269_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13269_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13269_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13274_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13274_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13274_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13274_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S14_13272_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S14_13272_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S14_13272_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S14_13272_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13274_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13274_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13274_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13274_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13274_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13274_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13274_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13274_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13279_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13279_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13279_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13279_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S15_13277_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S15_13277_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S15_13277_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S15_13277_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13279_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13279_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13279_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13279_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13279_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13279_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13279_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/SHL_u8_u8_13279_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13289_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13289_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13289_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13289_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13284_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13284_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13284_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13284_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S00_13282_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S00_13282_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S00_13282_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S00_13282_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13284_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13284_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13284_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13284_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13284_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13284_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13284_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13284_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13287_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13287_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13287_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13287_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S00x2_13285_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S00x2_13285_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S00x2_13285_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S00x2_13285_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13287_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13287_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13287_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13287_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13287_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13287_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13287_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13287_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S00x2_13288_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S06_13454_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S06_13454_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S06_13454_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13552_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S07_13455_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S07_13455_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S07_13455_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S07_13455_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13561_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13456_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13456_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13456_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13456_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13456_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13456_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S04_13322_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S04_13322_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S04_13322_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13324_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13324_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13324_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13324_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13324_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13324_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13324_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13324_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13327_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13327_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13327_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13327_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S04x2_13325_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S04x2_13325_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S04x2_13325_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S04x2_13325_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13327_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13327_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13327_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13327_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13327_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13327_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13327_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13327_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S04x2_13328_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S04x2_13328_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S04x2_13328_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S04x2_13328_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13329_start/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13329_start/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13329_start/req
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13329_start/ack
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13329_complete/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13329_complete/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13329_complete/req
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13329_complete/ack
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13339_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13339_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13339_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13339_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13334_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13334_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13334_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13334_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S05_13332_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S05_13332_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S05_13332_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S05_13332_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13334_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13334_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13334_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13334_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13334_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13334_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13334_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13334_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13337_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13337_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13337_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13337_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S05x2_13335_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S05x2_13335_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S05x2_13335_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S05x2_13335_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13337_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13337_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13337_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13337_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13337_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13337_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13337_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13337_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S05x2_13338_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S05x2_13338_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S05x2_13338_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S05x2_13338_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13339_start/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13339_start/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13339_start/req
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13339_start/ack
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13339_complete/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13339_complete/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13339_complete/req
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13339_complete/ack
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13349_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13349_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13349_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13349_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13344_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13344_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13344_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13344_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S06_13342_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S06_13342_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S06_13342_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S06_13342_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13344_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13344_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13344_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13344_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13344_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13344_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13344_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13344_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13347_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13347_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13347_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13347_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S06x2_13345_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S06x2_13345_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S06x2_13345_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S06x2_13345_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13347_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13347_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13347_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13347_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13347_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13347_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13347_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13347_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S06x2_13348_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S06x2_13348_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S06x2_13348_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S06x2_13348_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13349_start/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13349_start/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13349_start/req
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13349_start/ack
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13349_complete/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13349_complete/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13349_complete/req
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13349_complete/ack
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13359_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13359_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13359_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13359_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13354_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13354_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13354_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13354_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S07_13352_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S07_13352_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S07_13352_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S07_13352_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13354_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13354_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13354_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13354_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13354_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13354_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13354_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13354_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13357_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13357_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13357_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13357_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S07x2_13355_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S07x2_13355_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S07x2_13355_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S07x2_13355_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13357_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13357_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13357_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13357_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13357_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13357_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13357_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13357_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S07x2_13358_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S07x2_13358_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S07x2_13358_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S07x2_13358_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13359_start/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13359_start/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13359_start/req
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13359_start/ack
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13359_complete/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13359_complete/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13359_complete/req
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13359_complete/ack
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13369_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13369_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13369_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13369_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13364_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13364_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13364_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13364_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S08_13362_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S08_13362_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S08_13362_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S08_13362_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13364_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13364_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13364_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13364_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13364_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13364_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13364_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13364_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13367_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13367_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13367_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13367_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S08x2_13365_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S08x2_13365_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S08x2_13365_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S08x2_13365_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13448_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13564_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13367_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13367_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13444_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13367_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13367_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13367_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13367_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13444_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13367_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13367_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13447_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13453_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13447_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13448_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S08x2_13368_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S08x2_13368_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S08x2_13368_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S08x2_13368_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13447_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13447_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13369_start/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13369_start/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13444_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13369_start/req
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13369_start/ack
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13369_complete/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13369_complete/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13444_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13369_complete/req
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13369_complete/ack
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S03_13446_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S02_13445_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13379_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13379_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13379_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13379_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13374_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13374_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13374_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13374_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S09_13372_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S09_13372_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S09_13372_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S09_13372_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13447_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13564_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13447_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13374_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13374_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13448_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13374_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13374_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13374_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13374_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13448_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13374_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13374_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13444_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13444_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S04_13451_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S04_13451_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13444_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13457_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13377_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13377_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13377_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13377_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S09x2_13375_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S09x2_13375_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S09x2_13375_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S09x2_13375_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13447_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13377_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13377_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13448_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13377_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13377_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13377_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13377_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13448_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13377_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13377_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13444_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13453_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13444_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S09x2_13378_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S09x2_13378_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S09x2_13378_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S09x2_13378_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13447_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13564_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13447_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13447_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13379_start/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13379_start/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13439_complete/ack
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13379_start/req
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13379_start/ack
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13379_complete/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13379_complete/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13439_complete/req
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13379_complete/req
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13379_complete/ack
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S02_13445_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S02_13445_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13552_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13389_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13389_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13389_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13389_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13384_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13384_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13384_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13384_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S10_13382_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S10_13382_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S10_13382_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S10_13382_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13447_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Wc2_13562_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13444_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13384_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13384_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13439_complete/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13384_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13384_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13384_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13384_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13439_complete/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13384_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13384_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13444_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13444_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S05_13452_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S05_13452_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S01_13443_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13457_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13387_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13387_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13387_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13387_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S10x2_13385_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S10x2_13385_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S10x2_13385_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S10x2_13385_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13552_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13387_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13387_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13439_start/ack
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13387_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13387_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13387_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13387_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13439_start/req
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13387_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13387_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S01_13443_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13453_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S01_13443_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13552_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S10x2_13388_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S10x2_13388_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S10x2_13388_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S10x2_13388_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13669_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13389_start/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13389_start/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13439_start/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13389_start/req
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13389_start/ack
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13389_complete/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13389_complete/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13439_start/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13389_complete/req
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13389_complete/ack
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S02_13445_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13447_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13399_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13399_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13399_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13399_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13394_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13394_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13394_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13394_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S11_13392_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S11_13392_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S11_13392_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S11_13392_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13561_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13394_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13394_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13394_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13394_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13394_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13394_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13394_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13394_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Wc2_13553_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S09_13563_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S09_13563_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13552_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13555_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13565_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13397_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13397_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13397_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13397_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S11x2_13395_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S11x2_13395_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S11x2_13395_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S11x2_13395_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Wc2_13562_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13397_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13397_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13555_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13397_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13397_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13397_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13397_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13555_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13397_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13397_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13561_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13555_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S11x2_13398_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S11x2_13398_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S11x2_13398_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S11x2_13398_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S09x2g_13559_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13399_start/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13399_start/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13399_start/req
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13399_start/ack
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13399_complete/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13399_complete/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13399_complete/req
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13399_complete/ack
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13409_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13409_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13409_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13409_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13404_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13404_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13404_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13404_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S12_13402_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S12_13402_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S12_13402_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S12_13402_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Wc2_13562_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13552_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13561_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13404_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13404_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13404_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13404_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13404_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13404_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13404_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13404_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13561_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13565_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13561_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Wc2_13553_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13407_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13407_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13407_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13407_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S12x2_13405_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S12x2_13405_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S12x2_13405_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S12x2_13405_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Wc2_13553_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Wc2_13562_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S09_13563_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13561_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13407_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13407_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13556_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13407_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13407_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13407_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13407_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13407_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13407_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13564_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13564_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S09_13563_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S12x2_13408_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S12x2_13408_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S12x2_13408_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S12x2_13408_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13552_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13555_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13409_start/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13409_start/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13409_start/req
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13409_start/ack
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13409_complete/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13409_complete/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13409_complete/req
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13409_complete/ack
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13564_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13419_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13419_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13419_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13419_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13414_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13414_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13414_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13414_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S13_13412_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S13_13412_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S13_13412_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S13_13412_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13552_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13414_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13414_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13556_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13414_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13414_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13414_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13414_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13414_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13414_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13561_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13564_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13417_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13417_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13417_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13417_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S13x2_13415_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S13x2_13415_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S13x2_13415_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S13x2_13415_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13417_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13417_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13417_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13417_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13417_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13417_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13417_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13417_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S13x2_13418_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S13x2_13418_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S13x2_13418_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S13x2_13418_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13419_start/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13419_start/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13419_start/req
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13419_start/ack
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13419_complete/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13419_complete/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13419_complete/req
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13419_complete/ack
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13429_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13429_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13429_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13429_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13424_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13424_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13424_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13424_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S14_13422_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S14_13422_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S14_13422_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S14_13422_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13424_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13424_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13424_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13424_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13424_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13424_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13424_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13424_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13427_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13427_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13427_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13427_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S14x2_13425_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S14x2_13425_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S14x2_13425_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S14x2_13425_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13427_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13427_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13427_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13427_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13427_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13427_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13427_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13427_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S14x2_13428_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S14x2_13428_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S14x2_13428_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S14x2_13428_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13429_start/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13429_start/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13429_start/req
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13429_start/ack
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13429_complete/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13429_complete/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13429_complete/req
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13429_complete/ack
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13439_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13439_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13439_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13439_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13434_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13434_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13434_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13434_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S15_13432_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S15_13432_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S15_13432_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S15_13432_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13434_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13434_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13434_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13434_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13434_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13434_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13434_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/BITSEL_u8_u1_13434_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13437_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13437_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13437_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13437_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S15x2_13435_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S15x2_13435_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S15x2_13435_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S15x2_13435_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S05_13452_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S05_13452_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13453_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13453_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13453_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13453_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13453_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13453_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13453_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13453_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13456_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13456_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13456_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13456_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S06_13454_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13456_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13456_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13457_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13457_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13457_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13457_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13457_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13457_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13457_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13457_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13466_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13466_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13466_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13466_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13462_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13462_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13462_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13462_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S08_13460_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S08_13460_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S08_13460_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S08_13460_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S09_13461_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S09_13461_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S09_13461_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S09_13461_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13462_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13462_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13462_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13462_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13462_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13462_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13462_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13462_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13465_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13465_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13465_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13465_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S10_13463_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S10_13463_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S10_13463_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S10_13463_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S11_13464_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S11_13464_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S11_13464_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S11_13464_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13465_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13465_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13465_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13465_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13465_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13465_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13465_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13465_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13466_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13466_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13466_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13466_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13466_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13466_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13466_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13466_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13475_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13475_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13475_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13475_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13471_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13471_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13471_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13471_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S12_13469_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S12_13469_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S12_13469_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S12_13469_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S13_13470_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S13_13470_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S13_13470_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S13_13470_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13471_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13471_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13471_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13471_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13471_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13471_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13471_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13471_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13474_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13474_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13474_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13474_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S14_13472_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S14_13472_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S14_13472_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S14_13472_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S15_13473_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S15_13473_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S15_13473_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S15_13473_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13474_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13474_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13474_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13474_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13474_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13474_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13474_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13474_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13475_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13475_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13475_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13475_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13475_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13475_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13475_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13475_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13484_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13484_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13484_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13484_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13480_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13480_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13480_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13480_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S00x2g_13478_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S00x2g_13478_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S00x2g_13478_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S00x2g_13478_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S01x2g_13479_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S01x2g_13479_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S01x2g_13479_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S01x2g_13479_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13480_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13480_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13480_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13480_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13480_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13480_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13480_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13480_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13483_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13483_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13483_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13483_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Wc0_13481_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Wc0_13481_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Wc0_13481_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Wc0_13481_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S00_13482_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S00_13482_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S00_13482_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S00_13482_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13483_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13483_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13483_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13483_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13483_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13483_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13483_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13483_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13484_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13484_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13484_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13484_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13484_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13484_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13484_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13484_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13493_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13493_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13493_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13493_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13489_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13489_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13489_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13489_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S01x2g_13487_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S01x2g_13487_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S01x2g_13487_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S01x2g_13487_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S02x2g_13488_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S02x2g_13488_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S02x2g_13488_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S02x2g_13488_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13489_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13489_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13489_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13489_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13489_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13489_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13489_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13489_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13492_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13492_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13492_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13492_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Wc0_13490_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Wc0_13490_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Wc0_13490_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Wc0_13490_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S01_13491_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S01_13491_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S01_13491_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S01_13491_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13492_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13492_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13492_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13492_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13492_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13492_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13492_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13492_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13493_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13493_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13493_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13493_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13493_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13493_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13493_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13493_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13502_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13502_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13502_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13502_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13498_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13498_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13498_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13498_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S02x2g_13496_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S02x2g_13496_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S02x2g_13496_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S02x2g_13496_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S03x2g_13497_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S03x2g_13497_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S03x2g_13497_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S03x2g_13497_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13498_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13498_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13498_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13498_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13498_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13498_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13498_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13498_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13501_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13501_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13501_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13501_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Wc0_13499_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Wc0_13499_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Wc0_13499_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Wc0_13499_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13561_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S02_13500_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S02_13500_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S02_13500_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S02_13500_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13561_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_MX05_13677_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_MX06_13679_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13501_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13501_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13555_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13501_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13501_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13501_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13501_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13555_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13501_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13501_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13565_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13564_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13564_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13565_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13561_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S10x2g_13560_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13502_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13502_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13555_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13502_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13502_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13502_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13502_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13555_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13502_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13502_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13565_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13556_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S10x2g_13560_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13511_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13511_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13511_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13511_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13507_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13507_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13507_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13507_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S03x2g_13505_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S03x2g_13505_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S03x2g_13505_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S03x2g_13505_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Wc2_13553_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S10x2g_13560_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13556_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S00x2g_13506_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S00x2g_13506_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S00x2g_13506_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S00x2g_13506_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13555_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S10x2g_13560_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13556_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S09x2g_13559_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S09x2g_13559_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13507_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13507_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13555_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13507_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13507_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13507_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13507_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13555_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13507_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13507_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13556_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13564_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13556_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S09x2g_13559_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13510_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13510_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13510_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13510_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Wc0_13508_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Wc0_13508_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Wc0_13508_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Wc0_13508_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S03_13509_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S03_13509_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S03_13509_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S03_13509_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13669_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_MX04_13676_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13510_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13510_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S08_13554_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13510_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13510_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13510_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13510_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S08_13554_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13510_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13510_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13556_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13564_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13564_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13678_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13511_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13511_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S08_13554_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13511_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13511_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13511_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13511_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S08_13554_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13511_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13511_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13672_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13561_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13669_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13520_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13520_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13520_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13520_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13516_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13516_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13516_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13516_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S04x2g_13514_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S04x2g_13514_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S04x2g_13514_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S04x2g_13514_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_MX04_13676_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S05x2g_13515_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S05x2g_13515_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S05x2g_13515_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S05x2g_13515_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13516_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13516_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13516_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13516_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13516_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13516_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u16_u32_13673_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13516_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13516_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_MX06_13679_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_MX07_13680_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u16_u32_13682_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13678_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13519_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13519_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13519_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13519_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Wc1_13517_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Wc1_13517_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Wc1_13517_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Wc1_13517_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S04_13518_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S04_13518_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S04_13518_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S04_13518_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13672_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_MX03_13671_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13519_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13519_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13519_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13519_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13519_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13519_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13519_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13519_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13678_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13681_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13681_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13672_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13678_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13672_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13520_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13520_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13520_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13520_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13520_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13520_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13520_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13520_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_MX02_13670_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_MX04_13676_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13681_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13681_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_MX05_13677_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13529_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13529_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13529_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13529_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13525_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13525_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13525_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13525_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S05x2g_13523_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S05x2g_13523_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S05x2g_13523_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S05x2g_13523_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S06x2g_13524_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S06x2g_13524_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S06x2g_13524_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S06x2g_13524_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13672_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_MX07_13680_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13525_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13525_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u16_u32_13673_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13525_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13525_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13525_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13525_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13525_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13525_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13678_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13681_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13528_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13528_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13528_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13528_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Wc1_13526_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Wc1_13526_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Wc1_13526_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Wc1_13526_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_MX06_13679_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S05_13527_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S05_13527_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S05_13527_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S05_13527_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_MX07_13680_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_MX07_13680_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13672_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13528_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13528_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u16_u32_13673_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13528_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13528_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13528_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13528_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13528_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13528_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13669_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_MX03_13671_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_MX06_13679_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13529_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13529_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13529_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13529_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13529_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13529_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13669_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13529_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13529_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_MX03_13671_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13678_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_MX02_13670_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13538_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13538_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13538_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13538_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13534_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13534_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13534_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13534_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S06x2g_13532_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S06x2g_13532_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S06x2g_13532_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S06x2g_13532_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_MX03_13671_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13681_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13678_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S07x2g_13533_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S07x2g_13533_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S07x2g_13533_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S07x2g_13533_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13681_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_MX04_13676_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13672_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13534_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13534_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u16_u32_13673_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13534_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13534_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13534_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13534_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13534_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13534_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13681_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13537_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13537_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13537_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13537_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Wc1_13535_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Wc1_13535_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Wc1_13535_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Wc1_13535_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S06_13536_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S06_13536_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S06_13536_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S06_13536_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13537_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13537_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13537_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13537_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13537_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13537_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13537_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13537_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13538_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13538_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13538_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13538_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13538_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13538_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13538_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13538_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13547_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13547_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13547_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13547_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13543_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13543_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13543_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13543_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S07x2g_13541_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S07x2g_13541_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S07x2g_13541_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S07x2g_13541_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S04x2g_13542_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S04x2g_13542_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S04x2g_13542_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S04x2g_13542_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13543_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13543_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13543_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13543_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13543_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13543_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13543_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13543_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13546_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13546_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13546_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13546_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Wc1_13544_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Wc1_13544_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Wc1_13544_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Wc1_13544_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S07_13545_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S07_13545_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S07_13545_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S07_13545_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13546_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13546_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13546_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13546_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13546_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13546_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13546_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13546_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13547_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13547_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13547_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13547_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13547_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13547_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13547_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13547_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13556_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13556_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13556_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13556_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13552_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13552_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13552_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13552_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S08x2g_13550_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S08x2g_13550_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S08x2g_13550_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S08x2g_13550_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S09x2g_13551_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S09x2g_13551_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S09x2g_13551_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S09x2g_13551_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13565_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13565_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13565_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13565_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13565_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13565_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13565_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13574_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13574_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13574_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13574_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13570_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13570_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13570_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13570_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S10x2g_13568_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S10x2g_13568_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S10x2g_13568_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S10x2g_13568_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S11x2g_13569_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S11x2g_13569_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S11x2g_13569_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S11x2g_13569_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13570_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13570_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13570_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13570_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13570_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13570_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13570_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13570_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13573_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13573_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13573_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13573_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Wc2_13571_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Wc2_13571_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Wc2_13571_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Wc2_13571_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S10_13572_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S10_13572_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S10_13572_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S10_13572_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13573_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13573_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13573_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13573_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13573_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13573_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13573_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13573_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13574_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13574_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13574_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13574_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13574_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13574_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13574_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13574_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13583_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13583_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13583_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13583_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13579_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13579_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13579_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13579_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S11x2g_13577_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S11x2g_13577_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S11x2g_13577_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S11x2g_13577_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S08x2g_13578_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S08x2g_13578_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S08x2g_13578_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S08x2g_13578_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13579_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13579_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13579_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13579_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13579_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13579_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13579_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13579_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13582_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13582_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13582_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13582_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Wc2_13580_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Wc2_13580_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Wc2_13580_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Wc2_13580_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S11_13581_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S11_13581_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S11_13581_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S11_13581_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13582_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13582_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13582_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13582_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13582_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13582_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13582_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13582_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13583_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13583_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13583_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13583_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13583_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13583_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13583_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13583_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13592_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13592_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13592_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13592_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13588_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13588_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13588_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13588_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S12x2g_13586_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S12x2g_13586_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S12x2g_13586_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S12x2g_13586_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S13x2g_13587_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S13x2g_13587_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S13x2g_13587_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S13x2g_13587_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13588_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13588_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13588_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13588_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13588_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13588_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13588_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13588_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13591_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13591_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13591_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13591_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Wc3_13589_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Wc3_13589_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Wc3_13589_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Wc3_13589_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S12_13590_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S12_13590_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S12_13590_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S12_13590_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13591_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13591_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13591_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13591_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13591_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13591_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13591_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13591_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13592_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13592_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13592_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13592_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13592_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13592_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13592_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13592_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13601_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13601_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13601_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13601_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13597_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13597_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13597_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13597_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S13x2g_13595_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S13x2g_13595_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S13x2g_13595_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S13x2g_13595_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S14x2g_13596_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S14x2g_13596_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S14x2g_13596_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S14x2g_13596_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13597_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13597_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13597_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13597_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13597_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13597_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13597_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13597_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13600_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13600_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13600_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13600_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Wc3_13598_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Wc3_13598_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Wc3_13598_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Wc3_13598_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S13_13599_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S13_13599_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S13_13599_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S13_13599_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13600_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13600_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13600_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13600_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13600_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13600_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13600_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13600_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13601_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13601_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13601_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13601_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13601_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13601_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13601_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13601_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13610_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13610_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13610_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13610_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13606_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13606_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13606_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13606_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S14x2g_13604_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S14x2g_13604_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S14x2g_13604_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S14x2g_13604_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S15x2g_13605_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S15x2g_13605_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S15x2g_13605_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S15x2g_13605_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13606_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13606_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13606_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13606_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13606_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13606_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13606_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13606_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13609_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13609_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13609_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13609_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Wc3_13607_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Wc3_13607_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Wc3_13607_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Wc3_13607_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S14_13608_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S14_13608_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S14_13608_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S14_13608_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13609_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13609_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13609_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13609_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13609_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13609_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13609_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13609_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13610_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13610_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13610_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13610_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13610_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13610_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13610_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13610_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13619_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13619_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13619_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13619_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13615_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13615_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13615_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13615_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S15x2g_13613_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S15x2g_13613_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S15x2g_13613_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S15x2g_13613_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_MX02_13670_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13678_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u16_u32_13682_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S12x2g_13614_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S12x2g_13614_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S12x2g_13614_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S12x2g_13614_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_MX02_13670_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u16_u32_13682_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13678_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13678_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13615_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13615_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u16_u32_13673_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13615_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13615_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13615_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13615_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13672_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13615_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13615_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u16_u32_13682_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13681_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u16_u32_13673_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13678_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13618_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13618_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13618_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13618_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Wc3_13616_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Wc3_13616_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Wc3_13616_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Wc3_13616_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13678_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S15_13617_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S15_13617_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S15_13617_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S15_13617_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13618_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13618_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13672_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13618_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13618_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13618_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13618_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13672_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13618_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13618_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u16_u32_13673_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13681_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13681_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u16_u32_13673_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_MX05_13677_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_MX05_13677_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13619_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13619_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13672_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13619_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13619_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13619_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13619_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13672_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13619_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u8_u8_13619_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13681_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u16_u32_13628_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u16_u32_13628_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u16_u32_13628_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u16_u32_13628_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13624_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13624_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13624_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13624_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S00_13622_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S00_13622_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S00_13622_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S00_13622_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S01_13623_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S01_13623_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S01_13623_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S01_13623_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13624_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13624_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13624_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13624_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13624_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13624_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13624_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13624_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13627_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13627_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13627_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13627_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S02_13625_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S02_13625_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S02_13625_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S02_13625_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S03_13626_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S03_13626_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S03_13626_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S03_13626_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13627_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13627_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13627_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13627_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13627_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13627_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13627_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13627_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u16_u32_13628_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u16_u32_13628_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u16_u32_13628_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u16_u32_13628_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u16_u32_13628_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u16_u32_13628_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u16_u32_13628_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u16_u32_13628_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u16_u32_13637_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u16_u32_13637_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u16_u32_13637_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u16_u32_13637_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13633_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13633_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13633_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13633_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S04_13631_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S04_13631_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S04_13631_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S04_13631_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S05_13632_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S05_13632_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S05_13632_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S05_13632_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13633_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13633_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13633_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13633_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13633_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13633_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13633_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13633_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13636_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13636_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13636_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13636_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S06_13634_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S06_13634_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S06_13634_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S06_13634_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S07_13635_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S07_13635_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S07_13635_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S07_13635_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13636_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13636_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13636_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13636_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13636_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13636_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13636_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13636_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u16_u32_13637_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u16_u32_13637_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u16_u32_13637_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u16_u32_13637_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u16_u32_13637_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u16_u32_13637_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u16_u32_13637_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u16_u32_13637_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u16_u32_13646_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u16_u32_13646_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u16_u32_13646_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u16_u32_13646_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13642_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13642_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13642_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13642_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S08_13640_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S08_13640_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S08_13640_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S08_13640_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S09_13641_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S09_13641_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S09_13641_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S09_13641_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13642_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13642_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13642_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13642_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13642_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13642_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13642_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13642_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13645_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13645_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13645_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13645_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S10_13643_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S10_13643_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S10_13643_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S10_13643_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S11_13644_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S11_13644_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S11_13644_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S11_13644_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13645_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13645_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13645_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13645_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13645_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13645_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13645_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13645_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u16_u32_13646_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u16_u32_13646_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u16_u32_13646_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u16_u32_13646_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u16_u32_13646_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u16_u32_13646_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u16_u32_13646_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u16_u32_13646_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u16_u32_13655_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u16_u32_13655_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u16_u32_13655_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u16_u32_13655_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13651_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13651_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13651_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13651_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S12_13649_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S12_13649_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S12_13649_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S12_13649_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S13_13650_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S13_13650_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S13_13650_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S13_13650_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13651_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13651_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13651_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13651_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13651_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13651_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13651_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13651_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13654_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13654_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13654_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13654_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S14_13652_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S14_13652_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S14_13652_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S14_13652_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S15_13653_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S15_13653_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S15_13653_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_S15_13653_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13654_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13654_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13654_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13654_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13654_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13654_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13654_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13654_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u16_u32_13655_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u16_u32_13655_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u16_u32_13655_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u16_u32_13655_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u16_u32_13655_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u16_u32_13655_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u16_u32_13655_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u16_u32_13655_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u64_u128_13664_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u64_u128_13664_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u64_u128_13664_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u64_u128_13664_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u32_u64_13660_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u32_u64_13660_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u32_u64_13660_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u32_u64_13660_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Yl0_13658_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Yl0_13658_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Yl0_13658_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Yl0_13658_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Yl1_13659_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Yl1_13659_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Yl1_13659_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Yl1_13659_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u32_u64_13660_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u32_u64_13660_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u32_u64_13660_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u32_u64_13660_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u32_u64_13660_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u32_u64_13660_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u32_u64_13660_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u32_u64_13660_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u32_u64_13663_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u32_u64_13663_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u32_u64_13663_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u32_u64_13663_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Yl2_13661_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Yl2_13661_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Yl2_13661_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Yl2_13661_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Yl3_13662_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Yl3_13662_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Yl3_13662_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Yl3_13662_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u32_u64_13663_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u32_u64_13663_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u32_u64_13663_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u32_u64_13663_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u32_u64_13663_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u32_u64_13663_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u32_u64_13663_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u32_u64_13663_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u64_u128_13664_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u64_u128_13664_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u64_u128_13664_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u64_u128_13664_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u64_u128_13664_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u64_u128_13664_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u64_u128_13664_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u64_u128_13664_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u16_u32_13673_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u16_u32_13673_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u16_u32_13673_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u16_u32_13673_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13669_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13669_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13669_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13669_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_MX00_13667_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_MX00_13667_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_MX00_13667_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_MX00_13667_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_MX01_13668_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_MX01_13668_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_MX01_13668_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_MX01_13668_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13669_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13669_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13669_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u16_u32_13682_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u16_u32_13682_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u16_u32_13682_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u16_u32_13682_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u16_u32_13682_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u16_u32_13682_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u16_u32_13682_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u16_u32_13682_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u16_u32_13691_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u16_u32_13691_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u16_u32_13691_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u16_u32_13691_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13687_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13687_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13687_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13687_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_MX08_13685_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_MX08_13685_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_MX08_13685_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_MX08_13685_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_MX09_13686_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_MX09_13686_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_MX09_13686_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_MX09_13686_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13687_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13687_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13687_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13687_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13687_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13687_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13687_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13687_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13690_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13690_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13690_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13690_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_MX10_13688_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_MX10_13688_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_MX10_13688_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_MX10_13688_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_MX11_13689_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_MX11_13689_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_MX11_13689_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_MX11_13689_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13690_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13690_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13690_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13690_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13690_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13690_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13690_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13690_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u16_u32_13691_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u16_u32_13691_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u16_u32_13691_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u16_u32_13691_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u16_u32_13691_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u16_u32_13691_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u16_u32_13691_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u16_u32_13691_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u16_u32_13700_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u16_u32_13700_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u16_u32_13700_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u16_u32_13700_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13696_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13696_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13696_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13696_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_MX12_13694_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_MX12_13694_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_MX12_13694_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_MX12_13694_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_MX13_13695_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_MX13_13695_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_MX13_13695_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_MX13_13695_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13696_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13696_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13696_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13696_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13696_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13696_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13696_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13696_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13699_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13699_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13699_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13699_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_MX14_13697_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_MX14_13697_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_MX14_13697_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_MX14_13697_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_MX15_13698_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_MX15_13698_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_MX15_13698_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_MX15_13698_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13699_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13699_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13699_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13699_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13699_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13699_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13699_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u8_u16_13699_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u16_u32_13700_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u16_u32_13700_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u16_u32_13700_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u16_u32_13700_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u16_u32_13700_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u16_u32_13700_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u16_u32_13700_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u16_u32_13700_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u64_u128_13709_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u64_u128_13709_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u64_u128_13709_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u64_u128_13709_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u32_u64_13705_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u32_u64_13705_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u32_u64_13705_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u32_u64_13705_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Y0_13703_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Y0_13703_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Y0_13703_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Y0_13703_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Y1_13704_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Y1_13704_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Y1_13704_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Y1_13704_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u32_u64_13705_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u32_u64_13705_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u32_u64_13705_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u32_u64_13705_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u32_u64_13705_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u32_u64_13705_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u32_u64_13705_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u32_u64_13705_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u32_u64_13708_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u32_u64_13708_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u32_u64_13708_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u32_u64_13708_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Y2_13706_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Y2_13706_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Y2_13706_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Y2_13706_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Y3_13707_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Y3_13707_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Y3_13707_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Y3_13707_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u32_u64_13708_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u32_u64_13708_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u32_u64_13708_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u32_u64_13708_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u32_u64_13708_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u32_u64_13708_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u32_u64_13708_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u32_u64_13708_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u64_u128_13709_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u64_u128_13709_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u64_u128_13709_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u64_u128_13709_Sample/ra
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u64_u128_13709_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u64_u128_13709_Update/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u64_u128_13709_Update/cr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/CONCAT_u64_u128_13709_Update/ca
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13715_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13715_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13715_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13715_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_l_round_13712_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_l_round_13712_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_l_round_13712_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_l_round_13712_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Ylout_13713_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Ylout_13713_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Ylout_13713_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Ylout_13713_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Yout_13714_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Yout_13714_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Yout_13714_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Yout_13714_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13715_start/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13715_start/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13715_start/req
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13715_start/ack
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13715_complete/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13715_complete/$exit
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13715_complete/req
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/MUX_13715_complete/ack
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u128_u128_13720_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u128_u128_13720_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Zout_13718_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Zout_13718_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Zout_13718_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_Zout_13718_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_key_in_13719_sample_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_key_in_13719_sample_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_key_in_13719_update_start_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/R_key_in_13719_update_completed_
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u128_u128_13720_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u128_u128_13720_Sample/rr
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u128_u128_13720_Update/$entry
      -- CP-element group 0: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u128_u128_13720_Update/cr
      -- 
    cr_11103_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11103_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => enc_round_CP_7671_elements(0), ack => XOR_u128_u128_13720_inst_req_1); -- 
    rr_11098_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11098_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => enc_round_CP_7671_elements(0), ack => XOR_u128_u128_13720_inst_req_0); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u128_u128_13720_sample_completed_
      -- CP-element group 1: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u128_u128_13720_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u128_u128_13720_Sample/ra
      -- 
    ra_11099_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => XOR_u128_u128_13720_inst_ack_0, ack => enc_round_CP_7671_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2:  members (5) 
      -- CP-element group 2: 	 $exit
      -- CP-element group 2: 	 assign_stmt_13076_to_assign_stmt_13721/$exit
      -- CP-element group 2: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u128_u128_13720_update_completed_
      -- CP-element group 2: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u128_u128_13720_Update/$exit
      -- CP-element group 2: 	 assign_stmt_13076_to_assign_stmt_13721/XOR_u128_u128_13720_Update/ca
      -- 
    ca_11104_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => XOR_u128_u128_13720_inst_ack_1, ack => enc_round_CP_7671_elements(2)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal BITSEL_u8_u1_13284_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_13294_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_13304_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_13314_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_13324_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_13334_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_13344_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_13354_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_13364_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_13374_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_13384_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_13394_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_13404_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_13414_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_13424_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_13434_wire : std_logic_vector(0 downto 0);
    signal CONCAT_u32_u64_13660_wire : std_logic_vector(63 downto 0);
    signal CONCAT_u32_u64_13663_wire : std_logic_vector(63 downto 0);
    signal CONCAT_u32_u64_13705_wire : std_logic_vector(63 downto 0);
    signal CONCAT_u32_u64_13708_wire : std_logic_vector(63 downto 0);
    signal CONCAT_u8_u16_13624_wire : std_logic_vector(15 downto 0);
    signal CONCAT_u8_u16_13627_wire : std_logic_vector(15 downto 0);
    signal CONCAT_u8_u16_13633_wire : std_logic_vector(15 downto 0);
    signal CONCAT_u8_u16_13636_wire : std_logic_vector(15 downto 0);
    signal CONCAT_u8_u16_13642_wire : std_logic_vector(15 downto 0);
    signal CONCAT_u8_u16_13645_wire : std_logic_vector(15 downto 0);
    signal CONCAT_u8_u16_13651_wire : std_logic_vector(15 downto 0);
    signal CONCAT_u8_u16_13654_wire : std_logic_vector(15 downto 0);
    signal CONCAT_u8_u16_13669_wire : std_logic_vector(15 downto 0);
    signal CONCAT_u8_u16_13672_wire : std_logic_vector(15 downto 0);
    signal CONCAT_u8_u16_13678_wire : std_logic_vector(15 downto 0);
    signal CONCAT_u8_u16_13681_wire : std_logic_vector(15 downto 0);
    signal CONCAT_u8_u16_13687_wire : std_logic_vector(15 downto 0);
    signal CONCAT_u8_u16_13690_wire : std_logic_vector(15 downto 0);
    signal CONCAT_u8_u16_13696_wire : std_logic_vector(15 downto 0);
    signal CONCAT_u8_u16_13699_wire : std_logic_vector(15 downto 0);
    signal MX00_13485 : std_logic_vector(7 downto 0);
    signal MX01_13494 : std_logic_vector(7 downto 0);
    signal MX02_13503 : std_logic_vector(7 downto 0);
    signal MX03_13512 : std_logic_vector(7 downto 0);
    signal MX04_13521 : std_logic_vector(7 downto 0);
    signal MX05_13530 : std_logic_vector(7 downto 0);
    signal MX06_13539 : std_logic_vector(7 downto 0);
    signal MX07_13548 : std_logic_vector(7 downto 0);
    signal MX08_13557 : std_logic_vector(7 downto 0);
    signal MX09_13566 : std_logic_vector(7 downto 0);
    signal MX10_13575 : std_logic_vector(7 downto 0);
    signal MX11_13584 : std_logic_vector(7 downto 0);
    signal MX12_13593 : std_logic_vector(7 downto 0);
    signal MX13_13602 : std_logic_vector(7 downto 0);
    signal MX14_13611 : std_logic_vector(7 downto 0);
    signal MX15_13620 : std_logic_vector(7 downto 0);
    signal R_mod_const_13286_wire_constant : std_logic_vector(7 downto 0);
    signal R_mod_const_13296_wire_constant : std_logic_vector(7 downto 0);
    signal R_mod_const_13306_wire_constant : std_logic_vector(7 downto 0);
    signal R_mod_const_13316_wire_constant : std_logic_vector(7 downto 0);
    signal R_mod_const_13326_wire_constant : std_logic_vector(7 downto 0);
    signal R_mod_const_13336_wire_constant : std_logic_vector(7 downto 0);
    signal R_mod_const_13346_wire_constant : std_logic_vector(7 downto 0);
    signal R_mod_const_13356_wire_constant : std_logic_vector(7 downto 0);
    signal R_mod_const_13366_wire_constant : std_logic_vector(7 downto 0);
    signal R_mod_const_13376_wire_constant : std_logic_vector(7 downto 0);
    signal R_mod_const_13386_wire_constant : std_logic_vector(7 downto 0);
    signal R_mod_const_13396_wire_constant : std_logic_vector(7 downto 0);
    signal R_mod_const_13406_wire_constant : std_logic_vector(7 downto 0);
    signal R_mod_const_13416_wire_constant : std_logic_vector(7 downto 0);
    signal R_mod_const_13426_wire_constant : std_logic_vector(7 downto 0);
    signal R_mod_const_13436_wire_constant : std_logic_vector(7 downto 0);
    signal S00_13155 : std_logic_vector(7 downto 0);
    signal S00sr_13092 : std_logic_vector(7 downto 0);
    signal S00x2_13205 : std_logic_vector(7 downto 0);
    signal S00x2g_13290 : std_logic_vector(7 downto 0);
    signal S01_13158 : std_logic_vector(7 downto 0);
    signal S01sr_13096 : std_logic_vector(7 downto 0);
    signal S01x2_13210 : std_logic_vector(7 downto 0);
    signal S01x2g_13300 : std_logic_vector(7 downto 0);
    signal S02_13161 : std_logic_vector(7 downto 0);
    signal S02sr_13100 : std_logic_vector(7 downto 0);
    signal S02x2_13215 : std_logic_vector(7 downto 0);
    signal S02x2g_13310 : std_logic_vector(7 downto 0);
    signal S03_13164 : std_logic_vector(7 downto 0);
    signal S03sr_13104 : std_logic_vector(7 downto 0);
    signal S03x2_13220 : std_logic_vector(7 downto 0);
    signal S03x2g_13320 : std_logic_vector(7 downto 0);
    signal S04_13167 : std_logic_vector(7 downto 0);
    signal S04sr_13108 : std_logic_vector(7 downto 0);
    signal S04x2_13225 : std_logic_vector(7 downto 0);
    signal S04x2g_13330 : std_logic_vector(7 downto 0);
    signal S05_13170 : std_logic_vector(7 downto 0);
    signal S05sr_13112 : std_logic_vector(7 downto 0);
    signal S05x2_13230 : std_logic_vector(7 downto 0);
    signal S05x2g_13340 : std_logic_vector(7 downto 0);
    signal S06_13173 : std_logic_vector(7 downto 0);
    signal S06sr_13116 : std_logic_vector(7 downto 0);
    signal S06x2_13235 : std_logic_vector(7 downto 0);
    signal S06x2g_13350 : std_logic_vector(7 downto 0);
    signal S07_13176 : std_logic_vector(7 downto 0);
    signal S07sr_13120 : std_logic_vector(7 downto 0);
    signal S07x2_13240 : std_logic_vector(7 downto 0);
    signal S07x2g_13360 : std_logic_vector(7 downto 0);
    signal S08_13179 : std_logic_vector(7 downto 0);
    signal S08sr_13124 : std_logic_vector(7 downto 0);
    signal S08x2_13245 : std_logic_vector(7 downto 0);
    signal S08x2g_13370 : std_logic_vector(7 downto 0);
    signal S09_13182 : std_logic_vector(7 downto 0);
    signal S09sr_13128 : std_logic_vector(7 downto 0);
    signal S09x2_13250 : std_logic_vector(7 downto 0);
    signal S09x2g_13380 : std_logic_vector(7 downto 0);
    signal S10_13185 : std_logic_vector(7 downto 0);
    signal S10sr_13132 : std_logic_vector(7 downto 0);
    signal S10x2_13255 : std_logic_vector(7 downto 0);
    signal S10x2g_13390 : std_logic_vector(7 downto 0);
    signal S11_13188 : std_logic_vector(7 downto 0);
    signal S11sr_13136 : std_logic_vector(7 downto 0);
    signal S11x2_13260 : std_logic_vector(7 downto 0);
    signal S11x2g_13400 : std_logic_vector(7 downto 0);
    signal S12_13191 : std_logic_vector(7 downto 0);
    signal S12sr_13140 : std_logic_vector(7 downto 0);
    signal S12x2_13265 : std_logic_vector(7 downto 0);
    signal S12x2g_13410 : std_logic_vector(7 downto 0);
    signal S13_13194 : std_logic_vector(7 downto 0);
    signal S13sr_13144 : std_logic_vector(7 downto 0);
    signal S13x2_13270 : std_logic_vector(7 downto 0);
    signal S13x2g_13420 : std_logic_vector(7 downto 0);
    signal S14_13197 : std_logic_vector(7 downto 0);
    signal S14sr_13148 : std_logic_vector(7 downto 0);
    signal S14x2_13275 : std_logic_vector(7 downto 0);
    signal S14x2g_13430 : std_logic_vector(7 downto 0);
    signal S15_13200 : std_logic_vector(7 downto 0);
    signal S15sr_13152 : std_logic_vector(7 downto 0);
    signal S15x2_13280 : std_logic_vector(7 downto 0);
    signal S15x2g_13440 : std_logic_vector(7 downto 0);
    signal Sa_13076 : std_logic_vector(31 downto 0);
    signal Sb_13080 : std_logic_vector(31 downto 0);
    signal Sc_13084 : std_logic_vector(31 downto 0);
    signal Sd_13088 : std_logic_vector(31 downto 0);
    signal Wc0_13449 : std_logic_vector(7 downto 0);
    signal Wc1_13458 : std_logic_vector(7 downto 0);
    signal Wc2_13467 : std_logic_vector(7 downto 0);
    signal Wc3_13476 : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_13287_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_13297_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_13307_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_13317_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_13327_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_13337_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_13347_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_13357_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_13367_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_13377_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_13387_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_13397_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_13407_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_13417_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_13427_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_13437_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_13444_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_13447_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_13453_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_13456_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_13462_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_13465_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_13471_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_13474_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_13480_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_13483_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_13489_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_13492_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_13498_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_13501_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_13507_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_13510_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_13516_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_13519_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_13525_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_13528_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_13534_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_13537_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_13543_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_13546_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_13552_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_13555_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_13561_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_13564_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_13570_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_13573_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_13579_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_13582_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_13588_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_13591_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_13597_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_13600_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_13606_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_13609_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_13615_wire : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_13618_wire : std_logic_vector(7 downto 0);
    signal Y0_13674 : std_logic_vector(31 downto 0);
    signal Y1_13683 : std_logic_vector(31 downto 0);
    signal Y2_13692 : std_logic_vector(31 downto 0);
    signal Y3_13701 : std_logic_vector(31 downto 0);
    signal Yl0_13629 : std_logic_vector(31 downto 0);
    signal Yl1_13638 : std_logic_vector(31 downto 0);
    signal Yl2_13647 : std_logic_vector(31 downto 0);
    signal Yl3_13656 : std_logic_vector(31 downto 0);
    signal Ylout_13665 : std_logic_vector(127 downto 0);
    signal Yout_13710 : std_logic_vector(127 downto 0);
    signal Zout_13716 : std_logic_vector(127 downto 0);
    signal konst_13203_wire_constant : std_logic_vector(7 downto 0);
    signal konst_13208_wire_constant : std_logic_vector(7 downto 0);
    signal konst_13213_wire_constant : std_logic_vector(7 downto 0);
    signal konst_13218_wire_constant : std_logic_vector(7 downto 0);
    signal konst_13223_wire_constant : std_logic_vector(7 downto 0);
    signal konst_13228_wire_constant : std_logic_vector(7 downto 0);
    signal konst_13233_wire_constant : std_logic_vector(7 downto 0);
    signal konst_13238_wire_constant : std_logic_vector(7 downto 0);
    signal konst_13243_wire_constant : std_logic_vector(7 downto 0);
    signal konst_13248_wire_constant : std_logic_vector(7 downto 0);
    signal konst_13253_wire_constant : std_logic_vector(7 downto 0);
    signal konst_13258_wire_constant : std_logic_vector(7 downto 0);
    signal konst_13263_wire_constant : std_logic_vector(7 downto 0);
    signal konst_13268_wire_constant : std_logic_vector(7 downto 0);
    signal konst_13273_wire_constant : std_logic_vector(7 downto 0);
    signal konst_13278_wire_constant : std_logic_vector(7 downto 0);
    signal konst_13283_wire_constant : std_logic_vector(7 downto 0);
    signal konst_13293_wire_constant : std_logic_vector(7 downto 0);
    signal konst_13303_wire_constant : std_logic_vector(7 downto 0);
    signal konst_13313_wire_constant : std_logic_vector(7 downto 0);
    signal konst_13323_wire_constant : std_logic_vector(7 downto 0);
    signal konst_13333_wire_constant : std_logic_vector(7 downto 0);
    signal konst_13343_wire_constant : std_logic_vector(7 downto 0);
    signal konst_13353_wire_constant : std_logic_vector(7 downto 0);
    signal konst_13363_wire_constant : std_logic_vector(7 downto 0);
    signal konst_13373_wire_constant : std_logic_vector(7 downto 0);
    signal konst_13383_wire_constant : std_logic_vector(7 downto 0);
    signal konst_13393_wire_constant : std_logic_vector(7 downto 0);
    signal konst_13403_wire_constant : std_logic_vector(7 downto 0);
    signal konst_13413_wire_constant : std_logic_vector(7 downto 0);
    signal konst_13423_wire_constant : std_logic_vector(7 downto 0);
    signal konst_13433_wire_constant : std_logic_vector(7 downto 0);
    signal xxenc_roundxxmod_const : std_logic_vector(7 downto 0);
    signal xxenc_roundxxsel : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    R_mod_const_13286_wire_constant <= "00011011";
    R_mod_const_13296_wire_constant <= "00011011";
    R_mod_const_13306_wire_constant <= "00011011";
    R_mod_const_13316_wire_constant <= "00011011";
    R_mod_const_13326_wire_constant <= "00011011";
    R_mod_const_13336_wire_constant <= "00011011";
    R_mod_const_13346_wire_constant <= "00011011";
    R_mod_const_13356_wire_constant <= "00011011";
    R_mod_const_13366_wire_constant <= "00011011";
    R_mod_const_13376_wire_constant <= "00011011";
    R_mod_const_13386_wire_constant <= "00011011";
    R_mod_const_13396_wire_constant <= "00011011";
    R_mod_const_13406_wire_constant <= "00011011";
    R_mod_const_13416_wire_constant <= "00011011";
    R_mod_const_13426_wire_constant <= "00011011";
    R_mod_const_13436_wire_constant <= "00011011";
    konst_13203_wire_constant <= "00000001";
    konst_13208_wire_constant <= "00000001";
    konst_13213_wire_constant <= "00000001";
    konst_13218_wire_constant <= "00000001";
    konst_13223_wire_constant <= "00000001";
    konst_13228_wire_constant <= "00000001";
    konst_13233_wire_constant <= "00000001";
    konst_13238_wire_constant <= "00000001";
    konst_13243_wire_constant <= "00000001";
    konst_13248_wire_constant <= "00000001";
    konst_13253_wire_constant <= "00000001";
    konst_13258_wire_constant <= "00000001";
    konst_13263_wire_constant <= "00000001";
    konst_13268_wire_constant <= "00000001";
    konst_13273_wire_constant <= "00000001";
    konst_13278_wire_constant <= "00000001";
    konst_13283_wire_constant <= "00000111";
    konst_13293_wire_constant <= "00000111";
    konst_13303_wire_constant <= "00000111";
    konst_13313_wire_constant <= "00000111";
    konst_13323_wire_constant <= "00000111";
    konst_13333_wire_constant <= "00000111";
    konst_13343_wire_constant <= "00000111";
    konst_13353_wire_constant <= "00000111";
    konst_13363_wire_constant <= "00000111";
    konst_13373_wire_constant <= "00000111";
    konst_13383_wire_constant <= "00000111";
    konst_13393_wire_constant <= "00000111";
    konst_13403_wire_constant <= "00000111";
    konst_13413_wire_constant <= "00000111";
    konst_13423_wire_constant <= "00000111";
    konst_13433_wire_constant <= "00000111";
    xxenc_roundxxmod_const <= "00011011";
    xxenc_roundxxsel <= "01111111";
    -- flow-through select operator MUX_13289_inst
    S00x2g_13290 <= XOR_u8_u8_13287_wire when (BITSEL_u8_u1_13284_wire(0) /=  '0') else S00x2_13205;
    -- flow-through select operator MUX_13299_inst
    S01x2g_13300 <= XOR_u8_u8_13297_wire when (BITSEL_u8_u1_13294_wire(0) /=  '0') else S01x2_13210;
    -- flow-through select operator MUX_13309_inst
    S02x2g_13310 <= XOR_u8_u8_13307_wire when (BITSEL_u8_u1_13304_wire(0) /=  '0') else S02x2_13215;
    -- flow-through select operator MUX_13319_inst
    S03x2g_13320 <= XOR_u8_u8_13317_wire when (BITSEL_u8_u1_13314_wire(0) /=  '0') else S03x2_13220;
    -- flow-through select operator MUX_13329_inst
    S04x2g_13330 <= XOR_u8_u8_13327_wire when (BITSEL_u8_u1_13324_wire(0) /=  '0') else S04x2_13225;
    -- flow-through select operator MUX_13339_inst
    S05x2g_13340 <= XOR_u8_u8_13337_wire when (BITSEL_u8_u1_13334_wire(0) /=  '0') else S05x2_13230;
    -- flow-through select operator MUX_13349_inst
    S06x2g_13350 <= XOR_u8_u8_13347_wire when (BITSEL_u8_u1_13344_wire(0) /=  '0') else S06x2_13235;
    -- flow-through select operator MUX_13359_inst
    S07x2g_13360 <= XOR_u8_u8_13357_wire when (BITSEL_u8_u1_13354_wire(0) /=  '0') else S07x2_13240;
    -- flow-through select operator MUX_13369_inst
    S08x2g_13370 <= XOR_u8_u8_13367_wire when (BITSEL_u8_u1_13364_wire(0) /=  '0') else S08x2_13245;
    -- flow-through select operator MUX_13379_inst
    S09x2g_13380 <= XOR_u8_u8_13377_wire when (BITSEL_u8_u1_13374_wire(0) /=  '0') else S09x2_13250;
    -- flow-through select operator MUX_13389_inst
    S10x2g_13390 <= XOR_u8_u8_13387_wire when (BITSEL_u8_u1_13384_wire(0) /=  '0') else S10x2_13255;
    -- flow-through select operator MUX_13399_inst
    S11x2g_13400 <= XOR_u8_u8_13397_wire when (BITSEL_u8_u1_13394_wire(0) /=  '0') else S11x2_13260;
    -- flow-through select operator MUX_13409_inst
    S12x2g_13410 <= XOR_u8_u8_13407_wire when (BITSEL_u8_u1_13404_wire(0) /=  '0') else S12x2_13265;
    -- flow-through select operator MUX_13419_inst
    S13x2g_13420 <= XOR_u8_u8_13417_wire when (BITSEL_u8_u1_13414_wire(0) /=  '0') else S13x2_13270;
    -- flow-through select operator MUX_13429_inst
    S14x2g_13430 <= XOR_u8_u8_13427_wire when (BITSEL_u8_u1_13424_wire(0) /=  '0') else S14x2_13275;
    -- flow-through select operator MUX_13439_inst
    S15x2g_13440 <= XOR_u8_u8_13437_wire when (BITSEL_u8_u1_13434_wire(0) /=  '0') else S15x2_13280;
    -- flow-through select operator MUX_13715_inst
    Zout_13716 <= Ylout_13665 when (l_round_buffer(0) /=  '0') else Yout_13710;
    -- flow-through slice operator slice_13075_inst
    Sa_13076 <= round_in_buffer(127 downto 96);
    -- flow-through slice operator slice_13079_inst
    Sb_13080 <= round_in_buffer(95 downto 64);
    -- flow-through slice operator slice_13083_inst
    Sc_13084 <= round_in_buffer(63 downto 32);
    -- flow-through slice operator slice_13087_inst
    Sd_13088 <= round_in_buffer(31 downto 0);
    -- flow-through slice operator slice_13091_inst
    S00sr_13092 <= Sa_13076(31 downto 24);
    -- flow-through slice operator slice_13095_inst
    S01sr_13096 <= Sa_13076(23 downto 16);
    -- flow-through slice operator slice_13099_inst
    S02sr_13100 <= Sa_13076(15 downto 8);
    -- flow-through slice operator slice_13103_inst
    S03sr_13104 <= Sa_13076(7 downto 0);
    -- flow-through slice operator slice_13107_inst
    S04sr_13108 <= Sb_13080(31 downto 24);
    -- flow-through slice operator slice_13111_inst
    S05sr_13112 <= Sb_13080(23 downto 16);
    -- flow-through slice operator slice_13115_inst
    S06sr_13116 <= Sb_13080(15 downto 8);
    -- flow-through slice operator slice_13119_inst
    S07sr_13120 <= Sb_13080(7 downto 0);
    -- flow-through slice operator slice_13123_inst
    S08sr_13124 <= Sc_13084(31 downto 24);
    -- flow-through slice operator slice_13127_inst
    S09sr_13128 <= Sc_13084(23 downto 16);
    -- flow-through slice operator slice_13131_inst
    S10sr_13132 <= Sc_13084(15 downto 8);
    -- flow-through slice operator slice_13135_inst
    S11sr_13136 <= Sc_13084(7 downto 0);
    -- flow-through slice operator slice_13139_inst
    S12sr_13140 <= Sd_13088(31 downto 24);
    -- flow-through slice operator slice_13143_inst
    S13sr_13144 <= Sd_13088(23 downto 16);
    -- flow-through slice operator slice_13147_inst
    S14sr_13148 <= Sd_13088(15 downto 8);
    -- flow-through slice operator slice_13151_inst
    S15sr_13152 <= Sd_13088(7 downto 0);
    -- binary operator BITSEL_u8_u1_13284_inst
    process(S00_13155) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(S00_13155, konst_13283_wire_constant, tmp_var);
      BITSEL_u8_u1_13284_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_13294_inst
    process(S01_13158) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(S01_13158, konst_13293_wire_constant, tmp_var);
      BITSEL_u8_u1_13294_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_13304_inst
    process(S02_13161) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(S02_13161, konst_13303_wire_constant, tmp_var);
      BITSEL_u8_u1_13304_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_13314_inst
    process(S03_13164) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(S03_13164, konst_13313_wire_constant, tmp_var);
      BITSEL_u8_u1_13314_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_13324_inst
    process(S04_13167) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(S04_13167, konst_13323_wire_constant, tmp_var);
      BITSEL_u8_u1_13324_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_13334_inst
    process(S05_13170) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(S05_13170, konst_13333_wire_constant, tmp_var);
      BITSEL_u8_u1_13334_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_13344_inst
    process(S06_13173) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(S06_13173, konst_13343_wire_constant, tmp_var);
      BITSEL_u8_u1_13344_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_13354_inst
    process(S07_13176) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(S07_13176, konst_13353_wire_constant, tmp_var);
      BITSEL_u8_u1_13354_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_13364_inst
    process(S08_13179) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(S08_13179, konst_13363_wire_constant, tmp_var);
      BITSEL_u8_u1_13364_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_13374_inst
    process(S09_13182) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(S09_13182, konst_13373_wire_constant, tmp_var);
      BITSEL_u8_u1_13374_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_13384_inst
    process(S10_13185) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(S10_13185, konst_13383_wire_constant, tmp_var);
      BITSEL_u8_u1_13384_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_13394_inst
    process(S11_13188) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(S11_13188, konst_13393_wire_constant, tmp_var);
      BITSEL_u8_u1_13394_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_13404_inst
    process(S12_13191) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(S12_13191, konst_13403_wire_constant, tmp_var);
      BITSEL_u8_u1_13404_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_13414_inst
    process(S13_13194) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(S13_13194, konst_13413_wire_constant, tmp_var);
      BITSEL_u8_u1_13414_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_13424_inst
    process(S14_13197) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(S14_13197, konst_13423_wire_constant, tmp_var);
      BITSEL_u8_u1_13424_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_13434_inst
    process(S15_13200) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(S15_13200, konst_13433_wire_constant, tmp_var);
      BITSEL_u8_u1_13434_wire <= tmp_var; -- 
    end process;
    -- binary operator CONCAT_u16_u32_13628_inst
    process(CONCAT_u8_u16_13624_wire, CONCAT_u8_u16_13627_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u8_u16_13624_wire, CONCAT_u8_u16_13627_wire, tmp_var);
      Yl0_13629 <= tmp_var; -- 
    end process;
    -- binary operator CONCAT_u16_u32_13637_inst
    process(CONCAT_u8_u16_13633_wire, CONCAT_u8_u16_13636_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u8_u16_13633_wire, CONCAT_u8_u16_13636_wire, tmp_var);
      Yl1_13638 <= tmp_var; -- 
    end process;
    -- binary operator CONCAT_u16_u32_13646_inst
    process(CONCAT_u8_u16_13642_wire, CONCAT_u8_u16_13645_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u8_u16_13642_wire, CONCAT_u8_u16_13645_wire, tmp_var);
      Yl2_13647 <= tmp_var; -- 
    end process;
    -- binary operator CONCAT_u16_u32_13655_inst
    process(CONCAT_u8_u16_13651_wire, CONCAT_u8_u16_13654_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u8_u16_13651_wire, CONCAT_u8_u16_13654_wire, tmp_var);
      Yl3_13656 <= tmp_var; -- 
    end process;
    -- binary operator CONCAT_u16_u32_13673_inst
    process(CONCAT_u8_u16_13669_wire, CONCAT_u8_u16_13672_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u8_u16_13669_wire, CONCAT_u8_u16_13672_wire, tmp_var);
      Y0_13674 <= tmp_var; -- 
    end process;
    -- binary operator CONCAT_u16_u32_13682_inst
    process(CONCAT_u8_u16_13678_wire, CONCAT_u8_u16_13681_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u8_u16_13678_wire, CONCAT_u8_u16_13681_wire, tmp_var);
      Y1_13683 <= tmp_var; -- 
    end process;
    -- binary operator CONCAT_u16_u32_13691_inst
    process(CONCAT_u8_u16_13687_wire, CONCAT_u8_u16_13690_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u8_u16_13687_wire, CONCAT_u8_u16_13690_wire, tmp_var);
      Y2_13692 <= tmp_var; -- 
    end process;
    -- binary operator CONCAT_u16_u32_13700_inst
    process(CONCAT_u8_u16_13696_wire, CONCAT_u8_u16_13699_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u8_u16_13696_wire, CONCAT_u8_u16_13699_wire, tmp_var);
      Y3_13701 <= tmp_var; -- 
    end process;
    -- binary operator CONCAT_u32_u64_13660_inst
    process(Yl0_13629, Yl1_13638) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApConcat_proc(Yl0_13629, Yl1_13638, tmp_var);
      CONCAT_u32_u64_13660_wire <= tmp_var; -- 
    end process;
    -- binary operator CONCAT_u32_u64_13663_inst
    process(Yl2_13647, Yl3_13656) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApConcat_proc(Yl2_13647, Yl3_13656, tmp_var);
      CONCAT_u32_u64_13663_wire <= tmp_var; -- 
    end process;
    -- binary operator CONCAT_u32_u64_13705_inst
    process(Y0_13674, Y1_13683) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApConcat_proc(Y0_13674, Y1_13683, tmp_var);
      CONCAT_u32_u64_13705_wire <= tmp_var; -- 
    end process;
    -- binary operator CONCAT_u32_u64_13708_inst
    process(Y2_13692, Y3_13701) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApConcat_proc(Y2_13692, Y3_13701, tmp_var);
      CONCAT_u32_u64_13708_wire <= tmp_var; -- 
    end process;
    -- binary operator CONCAT_u64_u128_13664_inst
    process(CONCAT_u32_u64_13660_wire, CONCAT_u32_u64_13663_wire) -- 
      variable tmp_var : std_logic_vector(127 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u32_u64_13660_wire, CONCAT_u32_u64_13663_wire, tmp_var);
      Ylout_13665 <= tmp_var; -- 
    end process;
    -- binary operator CONCAT_u64_u128_13709_inst
    process(CONCAT_u32_u64_13705_wire, CONCAT_u32_u64_13708_wire) -- 
      variable tmp_var : std_logic_vector(127 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u32_u64_13705_wire, CONCAT_u32_u64_13708_wire, tmp_var);
      Yout_13710 <= tmp_var; -- 
    end process;
    -- binary operator CONCAT_u8_u16_13624_inst
    process(S00_13155, S01_13158) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApConcat_proc(S00_13155, S01_13158, tmp_var);
      CONCAT_u8_u16_13624_wire <= tmp_var; -- 
    end process;
    -- binary operator CONCAT_u8_u16_13627_inst
    process(S02_13161, S03_13164) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApConcat_proc(S02_13161, S03_13164, tmp_var);
      CONCAT_u8_u16_13627_wire <= tmp_var; -- 
    end process;
    -- binary operator CONCAT_u8_u16_13633_inst
    process(S04_13167, S05_13170) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApConcat_proc(S04_13167, S05_13170, tmp_var);
      CONCAT_u8_u16_13633_wire <= tmp_var; -- 
    end process;
    -- binary operator CONCAT_u8_u16_13636_inst
    process(S06_13173, S07_13176) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApConcat_proc(S06_13173, S07_13176, tmp_var);
      CONCAT_u8_u16_13636_wire <= tmp_var; -- 
    end process;
    -- binary operator CONCAT_u8_u16_13642_inst
    process(S08_13179, S09_13182) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApConcat_proc(S08_13179, S09_13182, tmp_var);
      CONCAT_u8_u16_13642_wire <= tmp_var; -- 
    end process;
    -- binary operator CONCAT_u8_u16_13645_inst
    process(S10_13185, S11_13188) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApConcat_proc(S10_13185, S11_13188, tmp_var);
      CONCAT_u8_u16_13645_wire <= tmp_var; -- 
    end process;
    -- binary operator CONCAT_u8_u16_13651_inst
    process(S12_13191, S13_13194) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApConcat_proc(S12_13191, S13_13194, tmp_var);
      CONCAT_u8_u16_13651_wire <= tmp_var; -- 
    end process;
    -- binary operator CONCAT_u8_u16_13654_inst
    process(S14_13197, S15_13200) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApConcat_proc(S14_13197, S15_13200, tmp_var);
      CONCAT_u8_u16_13654_wire <= tmp_var; -- 
    end process;
    -- binary operator CONCAT_u8_u16_13669_inst
    process(MX00_13485, MX01_13494) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApConcat_proc(MX00_13485, MX01_13494, tmp_var);
      CONCAT_u8_u16_13669_wire <= tmp_var; -- 
    end process;
    -- binary operator CONCAT_u8_u16_13672_inst
    process(MX02_13503, MX03_13512) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApConcat_proc(MX02_13503, MX03_13512, tmp_var);
      CONCAT_u8_u16_13672_wire <= tmp_var; -- 
    end process;
    -- binary operator CONCAT_u8_u16_13678_inst
    process(MX04_13521, MX05_13530) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApConcat_proc(MX04_13521, MX05_13530, tmp_var);
      CONCAT_u8_u16_13678_wire <= tmp_var; -- 
    end process;
    -- binary operator CONCAT_u8_u16_13681_inst
    process(MX06_13539, MX07_13548) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApConcat_proc(MX06_13539, MX07_13548, tmp_var);
      CONCAT_u8_u16_13681_wire <= tmp_var; -- 
    end process;
    -- binary operator CONCAT_u8_u16_13687_inst
    process(MX08_13557, MX09_13566) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApConcat_proc(MX08_13557, MX09_13566, tmp_var);
      CONCAT_u8_u16_13687_wire <= tmp_var; -- 
    end process;
    -- binary operator CONCAT_u8_u16_13690_inst
    process(MX10_13575, MX11_13584) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApConcat_proc(MX10_13575, MX11_13584, tmp_var);
      CONCAT_u8_u16_13690_wire <= tmp_var; -- 
    end process;
    -- binary operator CONCAT_u8_u16_13696_inst
    process(MX12_13593, MX13_13602) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApConcat_proc(MX12_13593, MX13_13602, tmp_var);
      CONCAT_u8_u16_13696_wire <= tmp_var; -- 
    end process;
    -- binary operator CONCAT_u8_u16_13699_inst
    process(MX14_13611, MX15_13620) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApConcat_proc(MX14_13611, MX15_13620, tmp_var);
      CONCAT_u8_u16_13699_wire <= tmp_var; -- 
    end process;
    -- binary operator SHL_u8_u8_13204_inst
    process(S00_13155) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntSHL_proc(S00_13155, konst_13203_wire_constant, tmp_var);
      S00x2_13205 <= tmp_var; -- 
    end process;
    -- binary operator SHL_u8_u8_13209_inst
    process(S01_13158) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntSHL_proc(S01_13158, konst_13208_wire_constant, tmp_var);
      S01x2_13210 <= tmp_var; -- 
    end process;
    -- binary operator SHL_u8_u8_13214_inst
    process(S02_13161) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntSHL_proc(S02_13161, konst_13213_wire_constant, tmp_var);
      S02x2_13215 <= tmp_var; -- 
    end process;
    -- binary operator SHL_u8_u8_13219_inst
    process(S03_13164) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntSHL_proc(S03_13164, konst_13218_wire_constant, tmp_var);
      S03x2_13220 <= tmp_var; -- 
    end process;
    -- binary operator SHL_u8_u8_13224_inst
    process(S04_13167) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntSHL_proc(S04_13167, konst_13223_wire_constant, tmp_var);
      S04x2_13225 <= tmp_var; -- 
    end process;
    -- binary operator SHL_u8_u8_13229_inst
    process(S05_13170) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntSHL_proc(S05_13170, konst_13228_wire_constant, tmp_var);
      S05x2_13230 <= tmp_var; -- 
    end process;
    -- binary operator SHL_u8_u8_13234_inst
    process(S06_13173) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntSHL_proc(S06_13173, konst_13233_wire_constant, tmp_var);
      S06x2_13235 <= tmp_var; -- 
    end process;
    -- binary operator SHL_u8_u8_13239_inst
    process(S07_13176) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntSHL_proc(S07_13176, konst_13238_wire_constant, tmp_var);
      S07x2_13240 <= tmp_var; -- 
    end process;
    -- binary operator SHL_u8_u8_13244_inst
    process(S08_13179) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntSHL_proc(S08_13179, konst_13243_wire_constant, tmp_var);
      S08x2_13245 <= tmp_var; -- 
    end process;
    -- binary operator SHL_u8_u8_13249_inst
    process(S09_13182) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntSHL_proc(S09_13182, konst_13248_wire_constant, tmp_var);
      S09x2_13250 <= tmp_var; -- 
    end process;
    -- binary operator SHL_u8_u8_13254_inst
    process(S10_13185) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntSHL_proc(S10_13185, konst_13253_wire_constant, tmp_var);
      S10x2_13255 <= tmp_var; -- 
    end process;
    -- binary operator SHL_u8_u8_13259_inst
    process(S11_13188) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntSHL_proc(S11_13188, konst_13258_wire_constant, tmp_var);
      S11x2_13260 <= tmp_var; -- 
    end process;
    -- binary operator SHL_u8_u8_13264_inst
    process(S12_13191) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntSHL_proc(S12_13191, konst_13263_wire_constant, tmp_var);
      S12x2_13265 <= tmp_var; -- 
    end process;
    -- binary operator SHL_u8_u8_13269_inst
    process(S13_13194) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntSHL_proc(S13_13194, konst_13268_wire_constant, tmp_var);
      S13x2_13270 <= tmp_var; -- 
    end process;
    -- binary operator SHL_u8_u8_13274_inst
    process(S14_13197) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntSHL_proc(S14_13197, konst_13273_wire_constant, tmp_var);
      S14x2_13275 <= tmp_var; -- 
    end process;
    -- binary operator SHL_u8_u8_13279_inst
    process(S15_13200) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntSHL_proc(S15_13200, konst_13278_wire_constant, tmp_var);
      S15x2_13280 <= tmp_var; -- 
    end process;
    -- shared split operator group (62) : XOR_u128_u128_13720_inst 
    ApIntXor_group_62: Block -- 
      signal data_in: std_logic_vector(255 downto 0);
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= Zout_13716 & key_in_buffer;
      round_out_buffer <= data_out(127 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= XOR_u128_u128_13720_inst_req_0;
      XOR_u128_u128_13720_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= XOR_u128_u128_13720_inst_req_1;
      XOR_u128_u128_13720_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(name => "gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntXor",
          name => "ApIntXor_group_62",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 128,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 128, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 128,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 62
    -- binary operator XOR_u8_u8_13287_inst
    process(S00x2_13205) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(S00x2_13205, R_mod_const_13286_wire_constant, tmp_var);
      XOR_u8_u8_13287_wire <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_13297_inst
    process(S01x2_13210) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(S01x2_13210, R_mod_const_13296_wire_constant, tmp_var);
      XOR_u8_u8_13297_wire <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_13307_inst
    process(S02x2_13215) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(S02x2_13215, R_mod_const_13306_wire_constant, tmp_var);
      XOR_u8_u8_13307_wire <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_13317_inst
    process(S03x2_13220) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(S03x2_13220, R_mod_const_13316_wire_constant, tmp_var);
      XOR_u8_u8_13317_wire <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_13327_inst
    process(S04x2_13225) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(S04x2_13225, R_mod_const_13326_wire_constant, tmp_var);
      XOR_u8_u8_13327_wire <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_13337_inst
    process(S05x2_13230) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(S05x2_13230, R_mod_const_13336_wire_constant, tmp_var);
      XOR_u8_u8_13337_wire <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_13347_inst
    process(S06x2_13235) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(S06x2_13235, R_mod_const_13346_wire_constant, tmp_var);
      XOR_u8_u8_13347_wire <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_13357_inst
    process(S07x2_13240) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(S07x2_13240, R_mod_const_13356_wire_constant, tmp_var);
      XOR_u8_u8_13357_wire <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_13367_inst
    process(S08x2_13245) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(S08x2_13245, R_mod_const_13366_wire_constant, tmp_var);
      XOR_u8_u8_13367_wire <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_13377_inst
    process(S09x2_13250) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(S09x2_13250, R_mod_const_13376_wire_constant, tmp_var);
      XOR_u8_u8_13377_wire <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_13387_inst
    process(S10x2_13255) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(S10x2_13255, R_mod_const_13386_wire_constant, tmp_var);
      XOR_u8_u8_13387_wire <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_13397_inst
    process(S11x2_13260) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(S11x2_13260, R_mod_const_13396_wire_constant, tmp_var);
      XOR_u8_u8_13397_wire <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_13407_inst
    process(S12x2_13265) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(S12x2_13265, R_mod_const_13406_wire_constant, tmp_var);
      XOR_u8_u8_13407_wire <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_13417_inst
    process(S13x2_13270) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(S13x2_13270, R_mod_const_13416_wire_constant, tmp_var);
      XOR_u8_u8_13417_wire <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_13427_inst
    process(S14x2_13275) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(S14x2_13275, R_mod_const_13426_wire_constant, tmp_var);
      XOR_u8_u8_13427_wire <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_13437_inst
    process(S15x2_13280) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(S15x2_13280, R_mod_const_13436_wire_constant, tmp_var);
      XOR_u8_u8_13437_wire <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_13444_inst
    process(S00_13155, S01_13158) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(S00_13155, S01_13158, tmp_var);
      XOR_u8_u8_13444_wire <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_13447_inst
    process(S02_13161, S03_13164) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(S02_13161, S03_13164, tmp_var);
      XOR_u8_u8_13447_wire <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_13448_inst
    process(XOR_u8_u8_13444_wire, XOR_u8_u8_13447_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(XOR_u8_u8_13444_wire, XOR_u8_u8_13447_wire, tmp_var);
      Wc0_13449 <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_13453_inst
    process(S04_13167, S05_13170) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(S04_13167, S05_13170, tmp_var);
      XOR_u8_u8_13453_wire <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_13456_inst
    process(S06_13173, S07_13176) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(S06_13173, S07_13176, tmp_var);
      XOR_u8_u8_13456_wire <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_13457_inst
    process(XOR_u8_u8_13453_wire, XOR_u8_u8_13456_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(XOR_u8_u8_13453_wire, XOR_u8_u8_13456_wire, tmp_var);
      Wc1_13458 <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_13462_inst
    process(S08_13179, S09_13182) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(S08_13179, S09_13182, tmp_var);
      XOR_u8_u8_13462_wire <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_13465_inst
    process(S10_13185, S11_13188) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(S10_13185, S11_13188, tmp_var);
      XOR_u8_u8_13465_wire <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_13466_inst
    process(XOR_u8_u8_13462_wire, XOR_u8_u8_13465_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(XOR_u8_u8_13462_wire, XOR_u8_u8_13465_wire, tmp_var);
      Wc2_13467 <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_13471_inst
    process(S12_13191, S13_13194) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(S12_13191, S13_13194, tmp_var);
      XOR_u8_u8_13471_wire <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_13474_inst
    process(S14_13197, S15_13200) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(S14_13197, S15_13200, tmp_var);
      XOR_u8_u8_13474_wire <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_13475_inst
    process(XOR_u8_u8_13471_wire, XOR_u8_u8_13474_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(XOR_u8_u8_13471_wire, XOR_u8_u8_13474_wire, tmp_var);
      Wc3_13476 <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_13480_inst
    process(S00x2g_13290, S01x2g_13300) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(S00x2g_13290, S01x2g_13300, tmp_var);
      XOR_u8_u8_13480_wire <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_13483_inst
    process(Wc0_13449, S00_13155) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(Wc0_13449, S00_13155, tmp_var);
      XOR_u8_u8_13483_wire <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_13484_inst
    process(XOR_u8_u8_13480_wire, XOR_u8_u8_13483_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(XOR_u8_u8_13480_wire, XOR_u8_u8_13483_wire, tmp_var);
      MX00_13485 <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_13489_inst
    process(S01x2g_13300, S02x2g_13310) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(S01x2g_13300, S02x2g_13310, tmp_var);
      XOR_u8_u8_13489_wire <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_13492_inst
    process(Wc0_13449, S01_13158) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(Wc0_13449, S01_13158, tmp_var);
      XOR_u8_u8_13492_wire <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_13493_inst
    process(XOR_u8_u8_13489_wire, XOR_u8_u8_13492_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(XOR_u8_u8_13489_wire, XOR_u8_u8_13492_wire, tmp_var);
      MX01_13494 <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_13498_inst
    process(S02x2g_13310, S03x2g_13320) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(S02x2g_13310, S03x2g_13320, tmp_var);
      XOR_u8_u8_13498_wire <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_13501_inst
    process(Wc0_13449, S02_13161) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(Wc0_13449, S02_13161, tmp_var);
      XOR_u8_u8_13501_wire <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_13502_inst
    process(XOR_u8_u8_13498_wire, XOR_u8_u8_13501_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(XOR_u8_u8_13498_wire, XOR_u8_u8_13501_wire, tmp_var);
      MX02_13503 <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_13507_inst
    process(S03x2g_13320, S00x2g_13290) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(S03x2g_13320, S00x2g_13290, tmp_var);
      XOR_u8_u8_13507_wire <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_13510_inst
    process(Wc0_13449, S03_13164) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(Wc0_13449, S03_13164, tmp_var);
      XOR_u8_u8_13510_wire <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_13511_inst
    process(XOR_u8_u8_13507_wire, XOR_u8_u8_13510_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(XOR_u8_u8_13507_wire, XOR_u8_u8_13510_wire, tmp_var);
      MX03_13512 <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_13516_inst
    process(S04x2g_13330, S05x2g_13340) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(S04x2g_13330, S05x2g_13340, tmp_var);
      XOR_u8_u8_13516_wire <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_13519_inst
    process(Wc1_13458, S04_13167) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(Wc1_13458, S04_13167, tmp_var);
      XOR_u8_u8_13519_wire <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_13520_inst
    process(XOR_u8_u8_13516_wire, XOR_u8_u8_13519_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(XOR_u8_u8_13516_wire, XOR_u8_u8_13519_wire, tmp_var);
      MX04_13521 <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_13525_inst
    process(S05x2g_13340, S06x2g_13350) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(S05x2g_13340, S06x2g_13350, tmp_var);
      XOR_u8_u8_13525_wire <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_13528_inst
    process(Wc1_13458, S05_13170) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(Wc1_13458, S05_13170, tmp_var);
      XOR_u8_u8_13528_wire <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_13529_inst
    process(XOR_u8_u8_13525_wire, XOR_u8_u8_13528_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(XOR_u8_u8_13525_wire, XOR_u8_u8_13528_wire, tmp_var);
      MX05_13530 <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_13534_inst
    process(S06x2g_13350, S07x2g_13360) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(S06x2g_13350, S07x2g_13360, tmp_var);
      XOR_u8_u8_13534_wire <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_13537_inst
    process(Wc1_13458, S06_13173) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(Wc1_13458, S06_13173, tmp_var);
      XOR_u8_u8_13537_wire <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_13538_inst
    process(XOR_u8_u8_13534_wire, XOR_u8_u8_13537_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(XOR_u8_u8_13534_wire, XOR_u8_u8_13537_wire, tmp_var);
      MX06_13539 <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_13543_inst
    process(S07x2g_13360, S04x2g_13330) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(S07x2g_13360, S04x2g_13330, tmp_var);
      XOR_u8_u8_13543_wire <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_13546_inst
    process(Wc1_13458, S07_13176) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(Wc1_13458, S07_13176, tmp_var);
      XOR_u8_u8_13546_wire <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_13547_inst
    process(XOR_u8_u8_13543_wire, XOR_u8_u8_13546_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(XOR_u8_u8_13543_wire, XOR_u8_u8_13546_wire, tmp_var);
      MX07_13548 <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_13552_inst
    process(S08x2g_13370, S09x2g_13380) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(S08x2g_13370, S09x2g_13380, tmp_var);
      XOR_u8_u8_13552_wire <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_13555_inst
    process(Wc2_13467, S08_13179) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(Wc2_13467, S08_13179, tmp_var);
      XOR_u8_u8_13555_wire <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_13556_inst
    process(XOR_u8_u8_13552_wire, XOR_u8_u8_13555_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(XOR_u8_u8_13552_wire, XOR_u8_u8_13555_wire, tmp_var);
      MX08_13557 <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_13561_inst
    process(S09x2g_13380, S10x2g_13390) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(S09x2g_13380, S10x2g_13390, tmp_var);
      XOR_u8_u8_13561_wire <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_13564_inst
    process(Wc2_13467, S09_13182) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(Wc2_13467, S09_13182, tmp_var);
      XOR_u8_u8_13564_wire <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_13565_inst
    process(XOR_u8_u8_13561_wire, XOR_u8_u8_13564_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(XOR_u8_u8_13561_wire, XOR_u8_u8_13564_wire, tmp_var);
      MX09_13566 <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_13570_inst
    process(S10x2g_13390, S11x2g_13400) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(S10x2g_13390, S11x2g_13400, tmp_var);
      XOR_u8_u8_13570_wire <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_13573_inst
    process(Wc2_13467, S10_13185) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(Wc2_13467, S10_13185, tmp_var);
      XOR_u8_u8_13573_wire <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_13574_inst
    process(XOR_u8_u8_13570_wire, XOR_u8_u8_13573_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(XOR_u8_u8_13570_wire, XOR_u8_u8_13573_wire, tmp_var);
      MX10_13575 <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_13579_inst
    process(S11x2g_13400, S08x2g_13370) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(S11x2g_13400, S08x2g_13370, tmp_var);
      XOR_u8_u8_13579_wire <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_13582_inst
    process(Wc2_13467, S11_13188) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(Wc2_13467, S11_13188, tmp_var);
      XOR_u8_u8_13582_wire <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_13583_inst
    process(XOR_u8_u8_13579_wire, XOR_u8_u8_13582_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(XOR_u8_u8_13579_wire, XOR_u8_u8_13582_wire, tmp_var);
      MX11_13584 <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_13588_inst
    process(S12x2g_13410, S13x2g_13420) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(S12x2g_13410, S13x2g_13420, tmp_var);
      XOR_u8_u8_13588_wire <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_13591_inst
    process(Wc3_13476, S12_13191) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(Wc3_13476, S12_13191, tmp_var);
      XOR_u8_u8_13591_wire <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_13592_inst
    process(XOR_u8_u8_13588_wire, XOR_u8_u8_13591_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(XOR_u8_u8_13588_wire, XOR_u8_u8_13591_wire, tmp_var);
      MX12_13593 <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_13597_inst
    process(S13x2g_13420, S14x2g_13430) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(S13x2g_13420, S14x2g_13430, tmp_var);
      XOR_u8_u8_13597_wire <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_13600_inst
    process(Wc3_13476, S13_13194) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(Wc3_13476, S13_13194, tmp_var);
      XOR_u8_u8_13600_wire <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_13601_inst
    process(XOR_u8_u8_13597_wire, XOR_u8_u8_13600_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(XOR_u8_u8_13597_wire, XOR_u8_u8_13600_wire, tmp_var);
      MX13_13602 <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_13606_inst
    process(S14x2g_13430, S15x2g_13440) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(S14x2g_13430, S15x2g_13440, tmp_var);
      XOR_u8_u8_13606_wire <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_13609_inst
    process(Wc3_13476, S14_13197) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(Wc3_13476, S14_13197, tmp_var);
      XOR_u8_u8_13609_wire <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_13610_inst
    process(XOR_u8_u8_13606_wire, XOR_u8_u8_13609_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(XOR_u8_u8_13606_wire, XOR_u8_u8_13609_wire, tmp_var);
      MX14_13611 <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_13615_inst
    process(S15x2g_13440, S12x2g_13410) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(S15x2g_13440, S12x2g_13410, tmp_var);
      XOR_u8_u8_13615_wire <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_13618_inst
    process(Wc3_13476, S15_13200) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(Wc3_13476, S15_13200, tmp_var);
      XOR_u8_u8_13618_wire <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_13619_inst
    process(XOR_u8_u8_13615_wire, XOR_u8_u8_13618_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(XOR_u8_u8_13615_wire, XOR_u8_u8_13618_wire, tmp_var);
      MX15_13620 <= tmp_var; -- 
    end process;
    call_inst_22628: sbox_mux_impl_Volatile port map(data_in => S00sr_13092, s_out => S00_13155); 
    call_inst_22629: sbox_mux_impl_Volatile port map(data_in => S05sr_13112, s_out => S01_13158); 
    call_inst_22630: sbox_mux_impl_Volatile port map(data_in => S10sr_13132, s_out => S02_13161); 
    call_inst_22631: sbox_mux_impl_Volatile port map(data_in => S15sr_13152, s_out => S03_13164); 
    call_inst_22632: sbox_mux_impl_Volatile port map(data_in => S04sr_13108, s_out => S04_13167); 
    call_inst_22633: sbox_mux_impl_Volatile port map(data_in => S09sr_13128, s_out => S05_13170); 
    call_inst_22634: sbox_mux_impl_Volatile port map(data_in => S14sr_13148, s_out => S06_13173); 
    call_inst_22635: sbox_mux_impl_Volatile port map(data_in => S03sr_13104, s_out => S07_13176); 
    call_inst_22636: sbox_mux_impl_Volatile port map(data_in => S08sr_13124, s_out => S08_13179); 
    call_inst_22637: sbox_mux_impl_Volatile port map(data_in => S13sr_13144, s_out => S09_13182); 
    call_inst_22638: sbox_mux_impl_Volatile port map(data_in => S02sr_13100, s_out => S10_13185); 
    call_inst_22639: sbox_mux_impl_Volatile port map(data_in => S07sr_13120, s_out => S11_13188); 
    call_inst_22640: sbox_mux_impl_Volatile port map(data_in => S12sr_13140, s_out => S12_13191); 
    call_inst_22641: sbox_mux_impl_Volatile port map(data_in => S01sr_13096, s_out => S13_13194); 
    call_inst_22642: sbox_mux_impl_Volatile port map(data_in => S06sr_13116, s_out => S14_13197); 
    call_inst_22643: sbox_mux_impl_Volatile port map(data_in => S11sr_13136, s_out => S15_13200); 
    -- 
  end Block; -- data_path
  -- 
end enc_round_Operator_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library work;
use work.ahir_system_global_package.all;
entity key_expand_single is -- 
  generic (tag_length : integer); 
  port ( -- 
    K_in : in  std_logic_vector(127 downto 0);
    Round_C : in  std_logic_vector(7 downto 0);
    K_out : out  std_logic_vector(127 downto 0);
    nRound_C : out  std_logic_vector(7 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity key_expand_single;
architecture key_expand_single_arch of key_expand_single is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 136)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 136)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal K_in_buffer :  std_logic_vector(127 downto 0);
  signal K_in_update_enable: Boolean;
  signal Round_C_buffer :  std_logic_vector(7 downto 0);
  signal Round_C_update_enable: Boolean;
  -- output port buffer signals
  signal K_out_buffer :  std_logic_vector(127 downto 0);
  signal K_out_update_enable: Boolean;
  signal nRound_C_buffer :  std_logic_vector(7 downto 0);
  signal nRound_C_update_enable: Boolean;
  signal key_expand_single_CP_2123_start: Boolean;
  signal key_expand_single_CP_2123_symbol: Boolean;
  -- volatile/operator module components. 
  component sbox_mux_impl_Volatile is -- 
    port ( -- 
      data_in : in  std_logic_vector(7 downto 0);
      s_out : out  std_logic_vector(7 downto 0)-- 
    );
    -- 
  end component; 
  -- links between control-path and data-path
  signal MUX_12146_inst_req_0 : boolean;
  signal MUX_12146_inst_ack_0 : boolean;
  signal MUX_12146_inst_req_1 : boolean;
  signal MUX_12146_inst_ack_1 : boolean;
  signal W_K_out_12148_inst_req_0 : boolean;
  signal W_K_out_12148_inst_ack_0 : boolean;
  signal W_K_out_12148_inst_req_1 : boolean;
  signal W_K_out_12148_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "key_expand_single_input_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      bypass_flag => true,
      data_width => tag_length + 136) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(127 downto 0) <= K_in;
  K_in_buffer <= in_buffer_data_out(127 downto 0);
  in_buffer_data_in(135 downto 128) <= Round_C;
  Round_C_buffer <= in_buffer_data_out(135 downto 128);
  in_buffer_data_in(tag_length + 135 downto 136) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 135 downto 136);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  key_expand_single_CP_2123_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "key_expand_single_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 136) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(127 downto 0) <= K_out_buffer;
  K_out <= out_buffer_data_out(127 downto 0);
  out_buffer_data_in(135 downto 128) <= nRound_C_buffer;
  nRound_C <= out_buffer_data_out(135 downto 128);
  out_buffer_data_in(tag_length + 135 downto 136) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 135 downto 136);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= key_expand_single_CP_2123_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= key_expand_single_CP_2123_start & tag_ilock_write_ack_symbol;
    gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= key_expand_single_CP_2123_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  key_expand_single_CP_2123: Block -- control-path 
    signal key_expand_single_CP_2123_elements: BooleanArray(5 downto 0);
    -- 
  begin -- 
    key_expand_single_CP_2123_elements(0) <= key_expand_single_CP_2123_start;
    key_expand_single_CP_2123_symbol <= key_expand_single_CP_2123_elements(5);
    -- CP-element group 0:  join  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	3 
    -- CP-element group 0: 	4 
    -- CP-element group 0:  members (1022) 
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11941_Update/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11913_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11913_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11925_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11925_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11921_Update/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11937_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K_in_11911_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11949_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_Ka_11932_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_Ka_11932_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11945_Update/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K12sr_12025_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11917_sample_completed_
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11945_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11937_Sample/rr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K_in_11911_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11917_Update/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11945_Update/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11913_Update/cr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K_in_11911_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11949_Update/cr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_Ka_11932_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11937_Update/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K12sr_12025_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11913_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11937_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11925_Update/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11913_Sample/rr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11929_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11949_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11913_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11913_Sample/ra
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11941_Update/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K_in_11911_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11937_Sample/ra
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11925_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_Ka_11932_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11913_Update/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11921_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_Kb_11944_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11913_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11933_Sample/ra
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11941_Update/ca
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11933_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11925_Sample/ra
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11921_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11925_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11925_Sample/rr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11925_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_Kb_11948_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11913_Update/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11949_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11933_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11949_Update/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_Ka_11928_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K_in_11924_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11917_Sample/ra
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK00_12030_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_Ka_11928_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11917_Sample/rr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11917_Update/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12016_Update/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11949_Update/ca
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11937_Update/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11917_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_Ka_11928_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11925_Update/cr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11921_Sample/ra
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_Kb_11944_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11917_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11913_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11933_Sample/rr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11917_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_Ka_11928_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11929_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11929_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11949_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11933_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11913_Update/ca
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11921_Sample/rr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K_in_11916_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11953_Sample/ra
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11929_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K_in_11916_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11941_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11953_Sample/rr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11949_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_Kb_11944_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K_in_11916_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12036_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11929_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K_in_11916_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_Kb_11944_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11917_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K_in_11924_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_Kb_11948_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11937_Update/ca
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11933_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11941_Update/cr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K_in_11924_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11937_Update/cr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11949_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11925_Update/ca
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_Kb_11952_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11917_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11925_Update/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K01_12014_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11925_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11945_Update/cr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11933_Update/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11921_Update/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12036_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11941_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11949_Sample/rr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11917_Update/cr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_Ka_11936_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11921_Update/cr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K03_12024_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11933_Update/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_Ka_11940_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_Ka_11940_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11921_Update/ca
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11953_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11933_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11933_Update/cr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11933_Update/ca
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_Kb_11948_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11941_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_Ka_11940_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11953_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_Ka_11940_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11929_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11917_Update/ca
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11921_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11945_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_Kb_11952_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11937_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11937_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11945_Update/ca
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_Ka_11936_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11941_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11945_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11929_Sample/rr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11945_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11945_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11929_Update/cr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK00_12030_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11953_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11921_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11953_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11921_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11945_Sample/rr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11929_Sample/ra
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12021_Update/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11929_Update/ca
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11941_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11933_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11937_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11953_Update/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11941_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11953_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11921_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11945_Sample/ra
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_Kb_11952_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K_in_11920_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11941_Sample/rr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11949_Sample/ra
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11937_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11949_Update/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12016_Update/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_Ka_11936_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_Kb_11952_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K_in_11924_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K_in_11920_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11929_Update/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11945_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K_in_11920_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K_in_11920_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11941_Sample/ra
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11929_Update/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11953_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K01_12014_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_Kb_11948_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_Ka_11936_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK06_12060_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K14sr_12015_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K03_12024_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12026_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K14sr_12015_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12061_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12061_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12031_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12016_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12016_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K14sr_12015_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K05_12034_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K12sr_12025_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_X0_12010_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12061_Sample/rr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12031_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12031_Update/cr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12016_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K05_12034_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K05_12034_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12011_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12031_Update/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12031_Sample/rr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12031_Update/ca
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12016_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K03_12024_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12011_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12011_Sample/rr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K05_12034_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK01_12035_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12016_Sample/rr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12016_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K03_12024_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12011_Sample/ra
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12021_Update/cr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12011_Update/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12031_Update/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK06_12060_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12011_Update/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K01_12014_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12016_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12021_Update/ca
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12026_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12056_Sample/rr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12026_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12061_Update/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12011_Update/cr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK06_12060_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12026_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K01_12014_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12016_Sample/ra
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12011_Update/ca
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12061_Sample/ra
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12026_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11953_Update/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11953_Update/cr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11953_Update/ca
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12056_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12056_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12066_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12066_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK05_12055_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11957_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11957_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11957_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11957_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_Kb_11956_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_Kb_11956_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_Kb_11956_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_Kb_11956_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK00_12030_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK05_12055_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK05_12055_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK05_12055_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K09_12054_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11957_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11957_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12021_Update/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11957_Sample/rr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11957_Sample/ra
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11957_Update/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11957_Update/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12021_Sample/ra
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11957_Update/cr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11957_Update/ca
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K09_12054_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K09_12054_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK07_12065_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK07_12065_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K09_12054_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12056_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11961_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11961_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11961_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11961_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_Kc_11960_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_Kc_11960_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_Kc_11960_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_Kc_11960_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK00_12030_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K10_12059_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12056_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12056_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12056_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11961_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11961_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12021_Sample/rr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11961_Sample/rr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11961_Sample/ra
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12066_Update/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12066_Update/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11961_Update/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11961_Update/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K14sr_12015_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11961_Update/cr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11961_Update/ca
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12051_Update/ca
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12051_Update/cr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK07_12065_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK07_12065_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12051_Update/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12051_Update/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11965_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11965_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11965_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11965_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_Kc_11964_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_Kc_11964_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_Kc_11964_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_Kc_11964_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K04_12029_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12051_Sample/ra
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12051_Sample/rr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12051_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11965_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11965_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12021_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11965_Sample/rr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11965_Sample/ra
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11965_Update/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11965_Update/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12021_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11965_Update/cr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11965_Update/ca
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12051_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K11_12064_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K11_12064_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK04_12050_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK04_12050_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11969_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11969_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11969_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11969_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_Kc_11968_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_Kc_11968_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_Kc_11968_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_Kc_11968_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K04_12029_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12036_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK04_12050_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK04_12050_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K08_12049_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11969_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11969_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K15sr_12020_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11969_Sample/rr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11969_Sample/ra
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11969_Update/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11969_Update/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K15sr_12020_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11969_Update/cr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11969_Update/ca
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K08_12049_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K08_12049_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K11_12064_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K11_12064_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K08_12049_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12051_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11973_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11973_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11973_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11973_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_Kc_11972_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_Kc_11972_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_Kc_11972_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_Kc_11972_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K04_12029_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12051_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12051_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12051_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12046_Update/ca
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11973_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11973_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K15sr_12020_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11973_Sample/rr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11973_Sample/ra
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11973_Update/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11973_Update/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K15sr_12020_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11973_Update/cr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11973_Update/ca
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12046_Update/cr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12046_Update/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12066_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12066_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12046_Update/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11977_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11977_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11977_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11977_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_Kd_11976_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_Kd_11976_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_Kd_11976_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_Kd_11976_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K04_12029_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K10_12059_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12046_Sample/ra
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12046_Sample/rr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12046_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11977_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11977_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K02_12019_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11977_Sample/rr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11977_Sample/ra
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11977_Update/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11977_Update/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K02_12019_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11977_Update/cr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11977_Update/ca
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12046_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12066_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12066_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK03_12045_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK03_12045_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11981_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11981_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11981_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11981_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_Kd_11980_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_Kd_11980_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_Kd_11980_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_Kd_11980_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12031_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK03_12045_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK03_12045_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K07_12044_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K07_12044_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11981_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11981_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K02_12019_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11981_Sample/rr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11981_Sample/ra
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11981_Update/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11981_Update/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K02_12019_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11981_Update/cr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11981_Update/ca
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K07_12044_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K07_12044_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12061_Update/ca
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12046_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12046_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11985_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11985_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11985_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11985_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_Kd_11984_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_Kd_11984_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_Kd_11984_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_Kd_11984_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12031_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12036_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12046_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12046_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12041_Update/ca
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11985_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11985_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12021_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11985_Sample/rr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11985_Sample/ra
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11985_Update/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11985_Update/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12021_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11985_Update/cr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11985_Update/ca
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12041_Update/cr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12041_Update/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12061_Update/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12061_Update/cr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12041_Update/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11989_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11989_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11989_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11989_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_Kd_11988_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_Kd_11988_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_Kd_11988_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_Kd_11988_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12031_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12041_Sample/ra
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12041_Sample/rr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12041_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12041_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11989_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11989_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12021_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11989_Sample/rr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11989_Sample/ra
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11989_Update/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11989_Update/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12021_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11989_Update/cr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/slice_11989_Update/ca
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK02_12040_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12066_Sample/rr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12066_Sample/ra
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK02_12040_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK02_12040_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/call_stmt_11993_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/call_stmt_11993_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/call_stmt_11993_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/call_stmt_11993_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12031_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K10_12059_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K10_12059_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K12_11991_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K12_11991_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K12_11991_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K12_11991_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12026_Update/ca
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK02_12040_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K06_12039_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K06_12039_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K06_12039_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/call_stmt_11996_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/call_stmt_11996_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/call_stmt_11996_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/call_stmt_11996_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12026_Update/cr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12061_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12061_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K13_11994_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K13_11994_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K13_11994_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K13_11994_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12026_Update/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K06_12039_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12041_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12041_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12041_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/call_stmt_11999_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/call_stmt_11999_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/call_stmt_11999_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/call_stmt_11999_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12026_Update/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12061_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12061_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K14_11997_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K14_11997_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K14_11997_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K14_11997_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12041_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12036_Update/ca
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12036_Update/cr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12036_Update/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/call_stmt_12002_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/call_stmt_12002_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/call_stmt_12002_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/call_stmt_12002_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12026_Sample/ra
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12056_Update/ca
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12056_Update/cr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K15_12000_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K15_12000_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K15_12000_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K15_12000_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12026_Sample/rr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12036_Update/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12036_Sample/ra
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12036_Sample/rr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12006_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12006_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12006_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12006_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_Round_C_12004_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_Round_C_12004_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_Round_C_12004_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_Round_C_12004_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K12sr_12025_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK01_12035_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12056_Update/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12056_Update/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K13sr_12005_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K13sr_12005_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K13sr_12005_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K13sr_12005_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12036_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12036_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK01_12035_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12006_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12006_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12016_Update/ca
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12006_Sample/rr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12006_Sample/ra
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12006_Update/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12006_Update/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12016_Update/cr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12006_Update/cr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12006_Update/ca
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK01_12035_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12056_Sample/ra
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK06_12060_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12026_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12031_Sample/ra
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12011_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12011_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12011_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12011_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K00_12009_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K00_12009_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K00_12009_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K00_12009_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_X0_12010_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_X0_12010_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_X0_12010_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK04_12098_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK04_12098_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK04_12098_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12066_Update/cr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12066_Update/ca
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12071_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12071_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12071_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12071_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K12_12069_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K12_12069_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K12_12069_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K12_12069_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK08_12070_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK08_12070_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK08_12070_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK08_12070_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12071_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12071_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12071_Sample/rr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12071_Sample/ra
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12071_Update/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12071_Update/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12071_Update/cr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12071_Update/ca
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12076_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12076_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12076_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12076_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K13_12074_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K13_12074_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K13_12074_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K13_12074_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK09_12075_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK09_12075_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK09_12075_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK09_12075_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12076_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12076_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12076_Sample/rr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12076_Sample/ra
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12076_Update/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12076_Update/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12076_Update/cr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12076_Update/ca
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12081_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12081_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12081_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12081_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K14_12079_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K14_12079_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K14_12079_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K14_12079_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK10_12080_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK10_12080_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK10_12080_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK10_12080_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12081_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12081_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12081_Sample/rr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12081_Sample/ra
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12081_Update/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12081_Update/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12081_Update/cr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12081_Update/ca
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12086_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12086_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12086_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12086_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K15_12084_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K15_12084_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K15_12084_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_K15_12084_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK11_12085_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK11_12085_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK11_12085_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK11_12085_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12086_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12086_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12086_Sample/rr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12086_Sample/ra
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12086_Update/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12086_Update/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12086_Update/cr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12086_Update/ca
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u16_u32_12095_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u16_u32_12095_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u16_u32_12095_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u16_u32_12095_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u8_u16_12091_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u8_u16_12091_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u8_u16_12091_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u8_u16_12091_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK00_12089_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK00_12089_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK00_12089_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK00_12089_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK01_12090_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK01_12090_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK01_12090_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK01_12090_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u8_u16_12091_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u8_u16_12091_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u8_u16_12091_Sample/rr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u8_u16_12091_Sample/ra
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u8_u16_12091_Update/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u8_u16_12091_Update/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u8_u16_12091_Update/cr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u8_u16_12091_Update/ca
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u8_u16_12094_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u8_u16_12094_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u8_u16_12094_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u8_u16_12094_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK02_12092_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK02_12092_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK02_12092_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK02_12092_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK03_12093_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK03_12093_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK03_12093_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK03_12093_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u8_u16_12094_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u8_u16_12094_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u8_u16_12094_Sample/rr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u8_u16_12094_Sample/ra
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u8_u16_12094_Update/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u8_u16_12094_Update/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u8_u16_12094_Update/cr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u8_u16_12094_Update/ca
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u16_u32_12095_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u16_u32_12095_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u16_u32_12095_Sample/rr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u16_u32_12095_Sample/ra
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u16_u32_12095_Update/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u16_u32_12095_Update/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u16_u32_12095_Update/cr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u16_u32_12095_Update/ca
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u16_u32_12104_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u16_u32_12104_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u16_u32_12104_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u16_u32_12104_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u8_u16_12100_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u8_u16_12100_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u8_u16_12100_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u8_u16_12100_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK04_12098_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK05_12099_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK05_12099_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK05_12099_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK05_12099_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u8_u16_12100_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u8_u16_12100_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u8_u16_12100_Sample/rr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u8_u16_12100_Sample/ra
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u8_u16_12100_Update/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u8_u16_12100_Update/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u8_u16_12100_Update/cr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u8_u16_12100_Update/ca
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u8_u16_12103_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u8_u16_12103_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u8_u16_12103_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u8_u16_12103_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK06_12101_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK06_12101_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK06_12101_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK06_12101_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK07_12102_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK07_12102_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK07_12102_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK07_12102_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u8_u16_12103_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u8_u16_12103_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u8_u16_12103_Sample/rr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u8_u16_12103_Sample/ra
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u8_u16_12103_Update/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u8_u16_12103_Update/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u8_u16_12103_Update/cr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u8_u16_12103_Update/ca
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u16_u32_12104_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u16_u32_12104_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u16_u32_12104_Sample/rr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u16_u32_12104_Sample/ra
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u16_u32_12104_Update/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u16_u32_12104_Update/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u16_u32_12104_Update/cr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u16_u32_12104_Update/ca
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u16_u32_12113_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u16_u32_12113_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u16_u32_12113_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u16_u32_12113_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u8_u16_12109_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u8_u16_12109_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u8_u16_12109_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u8_u16_12109_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK08_12107_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK08_12107_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK08_12107_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK08_12107_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK09_12108_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK09_12108_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK09_12108_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK09_12108_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u8_u16_12109_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u8_u16_12109_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u8_u16_12109_Sample/rr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u8_u16_12109_Sample/ra
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u8_u16_12109_Update/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u8_u16_12109_Update/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u8_u16_12109_Update/cr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u8_u16_12109_Update/ca
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u8_u16_12112_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u8_u16_12112_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u8_u16_12112_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u8_u16_12112_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK10_12110_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK10_12110_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK10_12110_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK10_12110_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK11_12111_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK11_12111_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK11_12111_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK11_12111_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u8_u16_12112_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u8_u16_12112_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u8_u16_12112_Sample/rr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u8_u16_12112_Sample/ra
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u8_u16_12112_Update/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u8_u16_12112_Update/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u8_u16_12112_Update/cr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u8_u16_12112_Update/ca
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u16_u32_12113_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u16_u32_12113_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u16_u32_12113_Sample/rr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u16_u32_12113_Sample/ra
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u16_u32_12113_Update/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u16_u32_12113_Update/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u16_u32_12113_Update/cr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u16_u32_12113_Update/ca
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u16_u32_12122_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u16_u32_12122_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u16_u32_12122_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u16_u32_12122_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u8_u16_12118_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u8_u16_12118_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u8_u16_12118_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u8_u16_12118_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK12_12116_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK12_12116_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK12_12116_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK12_12116_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK13_12117_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK13_12117_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK13_12117_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK13_12117_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u8_u16_12118_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u8_u16_12118_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u8_u16_12118_Sample/rr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u8_u16_12118_Sample/ra
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u8_u16_12118_Update/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u8_u16_12118_Update/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u8_u16_12118_Update/cr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u8_u16_12118_Update/ca
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u8_u16_12121_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u8_u16_12121_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u8_u16_12121_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u8_u16_12121_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK14_12119_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK14_12119_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK14_12119_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK14_12119_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK15_12120_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK15_12120_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK15_12120_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nK15_12120_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u8_u16_12121_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u8_u16_12121_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u8_u16_12121_Sample/rr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u8_u16_12121_Sample/ra
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u8_u16_12121_Update/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u8_u16_12121_Update/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u8_u16_12121_Update/cr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u8_u16_12121_Update/ca
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u16_u32_12122_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u16_u32_12122_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u16_u32_12122_Sample/rr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u16_u32_12122_Sample/ra
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u16_u32_12122_Update/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u16_u32_12122_Update/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u16_u32_12122_Update/cr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u16_u32_12122_Update/ca
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u64_u128_12131_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u64_u128_12131_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u64_u128_12131_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u64_u128_12131_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u32_u64_12127_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u32_u64_12127_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u32_u64_12127_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u32_u64_12127_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_Yk0_12125_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_Yk0_12125_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_Yk0_12125_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_Yk0_12125_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_Yk1_12126_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_Yk1_12126_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_Yk1_12126_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_Yk1_12126_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u32_u64_12127_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u32_u64_12127_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u32_u64_12127_Sample/rr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u32_u64_12127_Sample/ra
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u32_u64_12127_Update/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u32_u64_12127_Update/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u32_u64_12127_Update/cr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u32_u64_12127_Update/ca
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u32_u64_12130_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u32_u64_12130_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u32_u64_12130_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u32_u64_12130_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_Yk2_12128_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_Yk2_12128_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_Yk2_12128_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_Yk2_12128_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_Yk3_12129_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_Yk3_12129_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_Yk3_12129_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_Yk3_12129_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u32_u64_12130_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u32_u64_12130_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u32_u64_12130_Sample/rr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u32_u64_12130_Sample/ra
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u32_u64_12130_Update/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u32_u64_12130_Update/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u32_u64_12130_Update/cr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u32_u64_12130_Update/ca
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u64_u128_12131_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u64_u128_12131_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u64_u128_12131_Sample/rr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u64_u128_12131_Sample/ra
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u64_u128_12131_Update/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u64_u128_12131_Update/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u64_u128_12131_Update/cr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/CONCAT_u64_u128_12131_Update/ca
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/SHL_u8_u8_12136_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/SHL_u8_u8_12136_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/SHL_u8_u8_12136_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/SHL_u8_u8_12136_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_Round_C_12134_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_Round_C_12134_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_Round_C_12134_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_Round_C_12134_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/SHL_u8_u8_12136_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/SHL_u8_u8_12136_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/SHL_u8_u8_12136_Sample/rr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/SHL_u8_u8_12136_Sample/ra
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/SHL_u8_u8_12136_Update/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/SHL_u8_u8_12136_Update/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/SHL_u8_u8_12136_Update/cr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/SHL_u8_u8_12136_Update/ca
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/MUX_12146_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/MUX_12146_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/BITSEL_u8_u1_12141_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/BITSEL_u8_u1_12141_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/BITSEL_u8_u1_12141_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/BITSEL_u8_u1_12141_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_Round_C_12139_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_Round_C_12139_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_Round_C_12139_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_Round_C_12139_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/BITSEL_u8_u1_12141_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/BITSEL_u8_u1_12141_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/BITSEL_u8_u1_12141_Sample/rr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/BITSEL_u8_u1_12141_Sample/ra
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/BITSEL_u8_u1_12141_Update/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/BITSEL_u8_u1_12141_Update/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/BITSEL_u8_u1_12141_Update/cr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/BITSEL_u8_u1_12141_Update/ca
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12144_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12144_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12144_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12144_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_Rx2_12142_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_Rx2_12142_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_Rx2_12142_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_Rx2_12142_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12144_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12144_Sample/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12144_Sample/rr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12144_Sample/ra
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12144_Update/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12144_Update/$exit
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12144_Update/cr
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/XOR_u8_u8_12144_Update/ca
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_Rx2_12145_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_Rx2_12145_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_Rx2_12145_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_Rx2_12145_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/MUX_12146_start/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/MUX_12146_start/req
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/MUX_12146_complete/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/MUX_12146_complete/req
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nKey_12149_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nKey_12149_sample_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nKey_12149_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/R_nKey_12149_update_completed_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/assign_stmt_12150_sample_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/assign_stmt_12150_update_start_
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/assign_stmt_12150_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/assign_stmt_12150_Sample/req
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/assign_stmt_12150_Update/$entry
      -- CP-element group 0: 	 assign_stmt_11914_to_assign_stmt_12150/assign_stmt_12150_Update/req
      -- 
    req_3268_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3268_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => key_expand_single_CP_2123_elements(0), ack => W_K_out_12148_inst_req_0); -- 
    req_3255_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3255_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => key_expand_single_CP_2123_elements(0), ack => MUX_12146_inst_req_1); -- 
    req_3250_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3250_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => key_expand_single_CP_2123_elements(0), ack => MUX_12146_inst_req_0); -- 
    req_3273_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3273_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => key_expand_single_CP_2123_elements(0), ack => W_K_out_12148_inst_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 assign_stmt_11914_to_assign_stmt_12150/MUX_12146_sample_completed_
      -- CP-element group 1: 	 assign_stmt_11914_to_assign_stmt_12150/MUX_12146_start/$exit
      -- CP-element group 1: 	 assign_stmt_11914_to_assign_stmt_12150/MUX_12146_start/ack
      -- 
    ack_3251_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_12146_inst_ack_0, ack => key_expand_single_CP_2123_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	5 
    -- CP-element group 2:  members (3) 
      -- CP-element group 2: 	 assign_stmt_11914_to_assign_stmt_12150/MUX_12146_update_completed_
      -- CP-element group 2: 	 assign_stmt_11914_to_assign_stmt_12150/MUX_12146_complete/$exit
      -- CP-element group 2: 	 assign_stmt_11914_to_assign_stmt_12150/MUX_12146_complete/ack
      -- 
    ack_3256_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_12146_inst_ack_1, ack => key_expand_single_CP_2123_elements(2)); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	0 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 assign_stmt_11914_to_assign_stmt_12150/assign_stmt_12150_sample_completed_
      -- CP-element group 3: 	 assign_stmt_11914_to_assign_stmt_12150/assign_stmt_12150_Sample/$exit
      -- CP-element group 3: 	 assign_stmt_11914_to_assign_stmt_12150/assign_stmt_12150_Sample/ack
      -- 
    ack_3269_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_K_out_12148_inst_ack_0, ack => key_expand_single_CP_2123_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 assign_stmt_11914_to_assign_stmt_12150/assign_stmt_12150_update_completed_
      -- CP-element group 4: 	 assign_stmt_11914_to_assign_stmt_12150/assign_stmt_12150_Update/$exit
      -- CP-element group 4: 	 assign_stmt_11914_to_assign_stmt_12150/assign_stmt_12150_Update/ack
      -- 
    ack_3274_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_K_out_12148_inst_ack_1, ack => key_expand_single_CP_2123_elements(4)); -- 
    -- CP-element group 5:  join  transition  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	2 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (2) 
      -- CP-element group 5: 	 $exit
      -- CP-element group 5: 	 assign_stmt_11914_to_assign_stmt_12150/$exit
      -- 
    key_expand_single_cp_element_group_5: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 36) := "key_expand_single_cp_element_group_5"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= key_expand_single_CP_2123_elements(2) & key_expand_single_CP_2123_elements(4);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => key_expand_single_CP_2123_elements(5), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal BITSEL_u8_u1_12141_wire : std_logic_vector(0 downto 0);
    signal CONCAT_u32_u64_12127_wire : std_logic_vector(63 downto 0);
    signal CONCAT_u32_u64_12130_wire : std_logic_vector(63 downto 0);
    signal CONCAT_u8_u16_12091_wire : std_logic_vector(15 downto 0);
    signal CONCAT_u8_u16_12094_wire : std_logic_vector(15 downto 0);
    signal CONCAT_u8_u16_12100_wire : std_logic_vector(15 downto 0);
    signal CONCAT_u8_u16_12103_wire : std_logic_vector(15 downto 0);
    signal CONCAT_u8_u16_12109_wire : std_logic_vector(15 downto 0);
    signal CONCAT_u8_u16_12112_wire : std_logic_vector(15 downto 0);
    signal CONCAT_u8_u16_12118_wire : std_logic_vector(15 downto 0);
    signal CONCAT_u8_u16_12121_wire : std_logic_vector(15 downto 0);
    signal K00_11930 : std_logic_vector(7 downto 0);
    signal K01_11934 : std_logic_vector(7 downto 0);
    signal K02_11938 : std_logic_vector(7 downto 0);
    signal K03_11942 : std_logic_vector(7 downto 0);
    signal K04_11946 : std_logic_vector(7 downto 0);
    signal K05_11950 : std_logic_vector(7 downto 0);
    signal K06_11954 : std_logic_vector(7 downto 0);
    signal K07_11958 : std_logic_vector(7 downto 0);
    signal K08_11962 : std_logic_vector(7 downto 0);
    signal K09_11966 : std_logic_vector(7 downto 0);
    signal K10_11970 : std_logic_vector(7 downto 0);
    signal K11_11974 : std_logic_vector(7 downto 0);
    signal K12_11978 : std_logic_vector(7 downto 0);
    signal K12sr_11993 : std_logic_vector(7 downto 0);
    signal K13_11982 : std_logic_vector(7 downto 0);
    signal K13sr_11996 : std_logic_vector(7 downto 0);
    signal K14_11986 : std_logic_vector(7 downto 0);
    signal K14sr_11999 : std_logic_vector(7 downto 0);
    signal K15_11990 : std_logic_vector(7 downto 0);
    signal K15sr_12002 : std_logic_vector(7 downto 0);
    signal Ka_11914 : std_logic_vector(31 downto 0);
    signal Kb_11918 : std_logic_vector(31 downto 0);
    signal Kc_11922 : std_logic_vector(31 downto 0);
    signal Kd_11926 : std_logic_vector(31 downto 0);
    signal R_mod_const_12143_wire_constant : std_logic_vector(7 downto 0);
    signal Rx2_12137 : std_logic_vector(7 downto 0);
    signal X0_12007 : std_logic_vector(7 downto 0);
    signal XOR_u8_u8_12144_wire : std_logic_vector(7 downto 0);
    signal Yk0_12096 : std_logic_vector(31 downto 0);
    signal Yk1_12105 : std_logic_vector(31 downto 0);
    signal Yk2_12114 : std_logic_vector(31 downto 0);
    signal Yk3_12123 : std_logic_vector(31 downto 0);
    signal konst_12135_wire_constant : std_logic_vector(7 downto 0);
    signal konst_12140_wire_constant : std_logic_vector(7 downto 0);
    signal nK00_12012 : std_logic_vector(7 downto 0);
    signal nK01_12017 : std_logic_vector(7 downto 0);
    signal nK02_12022 : std_logic_vector(7 downto 0);
    signal nK03_12027 : std_logic_vector(7 downto 0);
    signal nK04_12032 : std_logic_vector(7 downto 0);
    signal nK05_12037 : std_logic_vector(7 downto 0);
    signal nK06_12042 : std_logic_vector(7 downto 0);
    signal nK07_12047 : std_logic_vector(7 downto 0);
    signal nK08_12052 : std_logic_vector(7 downto 0);
    signal nK09_12057 : std_logic_vector(7 downto 0);
    signal nK10_12062 : std_logic_vector(7 downto 0);
    signal nK11_12067 : std_logic_vector(7 downto 0);
    signal nK12_12072 : std_logic_vector(7 downto 0);
    signal nK13_12077 : std_logic_vector(7 downto 0);
    signal nK14_12082 : std_logic_vector(7 downto 0);
    signal nK15_12087 : std_logic_vector(7 downto 0);
    signal nKey_12132 : std_logic_vector(127 downto 0);
    signal xxkey_expand_singlexxmod_const : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    R_mod_const_12143_wire_constant <= "00011011";
    konst_12135_wire_constant <= "00000001";
    konst_12140_wire_constant <= "00000111";
    xxkey_expand_singlexxmod_const <= "00011011";
    MUX_12146_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= MUX_12146_inst_req_0;
      MUX_12146_inst_ack_0<= sample_ack(0);
      update_req(0) <= MUX_12146_inst_req_1;
      MUX_12146_inst_ack_1<= update_ack(0);
      MUX_12146_inst: SelectSplitProtocol generic map(name => "MUX_12146_inst", data_width => 8, buffering => 1, flow_through => false, full_rate => false) -- 
        port map( x => XOR_u8_u8_12144_wire, y => Rx2_12137, sel => BITSEL_u8_u1_12141_wire, z => nRound_C_buffer, sample_req => sample_req(0), sample_ack => sample_ack(0), update_req => update_req(0), update_ack => update_ack(0), clk => clk, reset => reset); -- 
      -- 
    end block;
    -- flow-through slice operator slice_11913_inst
    Ka_11914 <= K_in_buffer(127 downto 96);
    -- flow-through slice operator slice_11917_inst
    Kb_11918 <= K_in_buffer(95 downto 64);
    -- flow-through slice operator slice_11921_inst
    Kc_11922 <= K_in_buffer(63 downto 32);
    -- flow-through slice operator slice_11925_inst
    Kd_11926 <= K_in_buffer(31 downto 0);
    -- flow-through slice operator slice_11929_inst
    K00_11930 <= Ka_11914(31 downto 24);
    -- flow-through slice operator slice_11933_inst
    K01_11934 <= Ka_11914(23 downto 16);
    -- flow-through slice operator slice_11937_inst
    K02_11938 <= Ka_11914(15 downto 8);
    -- flow-through slice operator slice_11941_inst
    K03_11942 <= Ka_11914(7 downto 0);
    -- flow-through slice operator slice_11945_inst
    K04_11946 <= Kb_11918(31 downto 24);
    -- flow-through slice operator slice_11949_inst
    K05_11950 <= Kb_11918(23 downto 16);
    -- flow-through slice operator slice_11953_inst
    K06_11954 <= Kb_11918(15 downto 8);
    -- flow-through slice operator slice_11957_inst
    K07_11958 <= Kb_11918(7 downto 0);
    -- flow-through slice operator slice_11961_inst
    K08_11962 <= Kc_11922(31 downto 24);
    -- flow-through slice operator slice_11965_inst
    K09_11966 <= Kc_11922(23 downto 16);
    -- flow-through slice operator slice_11969_inst
    K10_11970 <= Kc_11922(15 downto 8);
    -- flow-through slice operator slice_11973_inst
    K11_11974 <= Kc_11922(7 downto 0);
    -- flow-through slice operator slice_11977_inst
    K12_11978 <= Kd_11926(31 downto 24);
    -- flow-through slice operator slice_11981_inst
    K13_11982 <= Kd_11926(23 downto 16);
    -- flow-through slice operator slice_11985_inst
    K14_11986 <= Kd_11926(15 downto 8);
    -- flow-through slice operator slice_11989_inst
    K15_11990 <= Kd_11926(7 downto 0);
    W_K_out_12148_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_K_out_12148_inst_req_0;
      W_K_out_12148_inst_ack_0<= wack(0);
      rreq(0) <= W_K_out_12148_inst_req_1;
      W_K_out_12148_inst_ack_1<= rack(0);
      W_K_out_12148_inst : InterlockBuffer generic map ( -- 
        name => "W_K_out_12148_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 128,
        out_data_width => 128,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nKey_12132,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => K_out_buffer,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- binary operator BITSEL_u8_u1_12141_inst
    process(Round_C_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(Round_C_buffer, konst_12140_wire_constant, tmp_var);
      BITSEL_u8_u1_12141_wire <= tmp_var; -- 
    end process;
    -- binary operator CONCAT_u16_u32_12095_inst
    process(CONCAT_u8_u16_12091_wire, CONCAT_u8_u16_12094_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u8_u16_12091_wire, CONCAT_u8_u16_12094_wire, tmp_var);
      Yk0_12096 <= tmp_var; -- 
    end process;
    -- binary operator CONCAT_u16_u32_12104_inst
    process(CONCAT_u8_u16_12100_wire, CONCAT_u8_u16_12103_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u8_u16_12100_wire, CONCAT_u8_u16_12103_wire, tmp_var);
      Yk1_12105 <= tmp_var; -- 
    end process;
    -- binary operator CONCAT_u16_u32_12113_inst
    process(CONCAT_u8_u16_12109_wire, CONCAT_u8_u16_12112_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u8_u16_12109_wire, CONCAT_u8_u16_12112_wire, tmp_var);
      Yk2_12114 <= tmp_var; -- 
    end process;
    -- binary operator CONCAT_u16_u32_12122_inst
    process(CONCAT_u8_u16_12118_wire, CONCAT_u8_u16_12121_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u8_u16_12118_wire, CONCAT_u8_u16_12121_wire, tmp_var);
      Yk3_12123 <= tmp_var; -- 
    end process;
    -- binary operator CONCAT_u32_u64_12127_inst
    process(Yk0_12096, Yk1_12105) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApConcat_proc(Yk0_12096, Yk1_12105, tmp_var);
      CONCAT_u32_u64_12127_wire <= tmp_var; -- 
    end process;
    -- binary operator CONCAT_u32_u64_12130_inst
    process(Yk2_12114, Yk3_12123) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApConcat_proc(Yk2_12114, Yk3_12123, tmp_var);
      CONCAT_u32_u64_12130_wire <= tmp_var; -- 
    end process;
    -- binary operator CONCAT_u64_u128_12131_inst
    process(CONCAT_u32_u64_12127_wire, CONCAT_u32_u64_12130_wire) -- 
      variable tmp_var : std_logic_vector(127 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u32_u64_12127_wire, CONCAT_u32_u64_12130_wire, tmp_var);
      nKey_12132 <= tmp_var; -- 
    end process;
    -- binary operator CONCAT_u8_u16_12091_inst
    process(nK00_12012, nK01_12017) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApConcat_proc(nK00_12012, nK01_12017, tmp_var);
      CONCAT_u8_u16_12091_wire <= tmp_var; -- 
    end process;
    -- binary operator CONCAT_u8_u16_12094_inst
    process(nK02_12022, nK03_12027) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApConcat_proc(nK02_12022, nK03_12027, tmp_var);
      CONCAT_u8_u16_12094_wire <= tmp_var; -- 
    end process;
    -- binary operator CONCAT_u8_u16_12100_inst
    process(nK04_12032, nK05_12037) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApConcat_proc(nK04_12032, nK05_12037, tmp_var);
      CONCAT_u8_u16_12100_wire <= tmp_var; -- 
    end process;
    -- binary operator CONCAT_u8_u16_12103_inst
    process(nK06_12042, nK07_12047) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApConcat_proc(nK06_12042, nK07_12047, tmp_var);
      CONCAT_u8_u16_12103_wire <= tmp_var; -- 
    end process;
    -- binary operator CONCAT_u8_u16_12109_inst
    process(nK08_12052, nK09_12057) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApConcat_proc(nK08_12052, nK09_12057, tmp_var);
      CONCAT_u8_u16_12109_wire <= tmp_var; -- 
    end process;
    -- binary operator CONCAT_u8_u16_12112_inst
    process(nK10_12062, nK11_12067) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApConcat_proc(nK10_12062, nK11_12067, tmp_var);
      CONCAT_u8_u16_12112_wire <= tmp_var; -- 
    end process;
    -- binary operator CONCAT_u8_u16_12118_inst
    process(nK12_12072, nK13_12077) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApConcat_proc(nK12_12072, nK13_12077, tmp_var);
      CONCAT_u8_u16_12118_wire <= tmp_var; -- 
    end process;
    -- binary operator CONCAT_u8_u16_12121_inst
    process(nK14_12082, nK15_12087) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApConcat_proc(nK14_12082, nK15_12087, tmp_var);
      CONCAT_u8_u16_12121_wire <= tmp_var; -- 
    end process;
    -- binary operator SHL_u8_u8_12136_inst
    process(Round_C_buffer) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntSHL_proc(Round_C_buffer, konst_12135_wire_constant, tmp_var);
      Rx2_12137 <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_12006_inst
    process(Round_C_buffer, K13sr_11996) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(Round_C_buffer, K13sr_11996, tmp_var);
      X0_12007 <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_12011_inst
    process(K00_11930, X0_12007) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(K00_11930, X0_12007, tmp_var);
      nK00_12012 <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_12016_inst
    process(K01_11934, K14sr_11999) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(K01_11934, K14sr_11999, tmp_var);
      nK01_12017 <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_12021_inst
    process(K02_11938, K15sr_12002) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(K02_11938, K15sr_12002, tmp_var);
      nK02_12022 <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_12026_inst
    process(K03_11942, K12sr_11993) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(K03_11942, K12sr_11993, tmp_var);
      nK03_12027 <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_12031_inst
    process(K04_11946, nK00_12012) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(K04_11946, nK00_12012, tmp_var);
      nK04_12032 <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_12036_inst
    process(K05_11950, nK01_12017) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(K05_11950, nK01_12017, tmp_var);
      nK05_12037 <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_12041_inst
    process(K06_11954, nK02_12022) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(K06_11954, nK02_12022, tmp_var);
      nK06_12042 <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_12046_inst
    process(K07_11958, nK03_12027) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(K07_11958, nK03_12027, tmp_var);
      nK07_12047 <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_12051_inst
    process(K08_11962, nK04_12032) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(K08_11962, nK04_12032, tmp_var);
      nK08_12052 <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_12056_inst
    process(K09_11966, nK05_12037) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(K09_11966, nK05_12037, tmp_var);
      nK09_12057 <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_12061_inst
    process(K10_11970, nK06_12042) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(K10_11970, nK06_12042, tmp_var);
      nK10_12062 <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_12066_inst
    process(K11_11974, nK07_12047) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(K11_11974, nK07_12047, tmp_var);
      nK11_12067 <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_12071_inst
    process(K12_11978, nK08_12052) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(K12_11978, nK08_12052, tmp_var);
      nK12_12072 <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_12076_inst
    process(K13_11982, nK09_12057) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(K13_11982, nK09_12057, tmp_var);
      nK13_12077 <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_12081_inst
    process(K14_11986, nK10_12062) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(K14_11986, nK10_12062, tmp_var);
      nK14_12082 <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_12086_inst
    process(K15_11990, nK11_12067) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(K15_11990, nK11_12067, tmp_var);
      nK15_12087 <= tmp_var; -- 
    end process;
    -- binary operator XOR_u8_u8_12144_inst
    process(Rx2_12137) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntXor_proc(Rx2_12137, R_mod_const_12143_wire_constant, tmp_var);
      XOR_u8_u8_12144_wire <= tmp_var; -- 
    end process;
    call_inst_13901: sbox_mux_impl_Volatile port map(data_in => K12_11978, s_out => K12sr_11993); 
    call_inst_13902: sbox_mux_impl_Volatile port map(data_in => K13_11982, s_out => K13sr_11996); 
    call_inst_13903: sbox_mux_impl_Volatile port map(data_in => K14_11986, s_out => K14sr_11999); 
    call_inst_13904: sbox_mux_impl_Volatile port map(data_in => K15_11990, s_out => K15sr_12002); 
    -- 
  end Block; -- data_path
  -- 
end key_expand_single_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library work;
use work.ahir_system_global_package.all;
entity sbox_mux_impl_Volatile is -- 
  port ( -- 
    data_in : in  std_logic_vector(7 downto 0);
    s_out : out  std_logic_vector(7 downto 0)-- 
  );
  -- 
end entity sbox_mux_impl_Volatile;
architecture sbox_mux_impl_Volatile_arch of sbox_mux_impl_Volatile is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector(8-1 downto 0);
  signal default_zero_sig: std_logic;
  -- input port buffer signals
  signal data_in_buffer :  std_logic_vector(7 downto 0);
  -- output port buffer signals
  signal s_out_buffer :  std_logic_vector(7 downto 0);
  -- volatile/operator module components. 
  -- 
begin --  
  -- input handling ------------------------------------------------
  data_in_buffer <= data_in;
  -- output handling  -------------------------------------------------------
  s_out <= s_out_buffer;
  -- the control path --------------------------------------------------
  default_zero_sig <= '0';
  -- volatile module, no control path
  -- the data path
  data_path: Block -- 
    signal BITSEL_u8_u1_10008_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_10018_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_10028_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_10038_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_10048_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_10058_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_10068_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_10078_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_10088_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_10098_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_10108_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_10118_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_10128_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_10138_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_10148_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_10158_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_10168_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_10178_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_10188_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_10198_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_10208_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_10218_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_10228_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_10238_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_10248_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_10258_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_10268_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_10278_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_10288_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_10298_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_10308_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_10318_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_10328_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_10338_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_10348_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_10358_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_10368_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_10378_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_10388_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_10398_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_10408_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_10418_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_10428_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_10438_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_10448_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_10458_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_10468_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_10478_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_10488_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_10498_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_10508_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_10518_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_10528_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_10538_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_10548_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_10558_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_10568_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_10578_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_10588_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_10598_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_10608_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_10618_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_10628_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_10638_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_10648_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_10658_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_10668_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_10678_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_10688_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_10698_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_10708_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_10718_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_10728_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_10738_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_10748_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_10758_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_10768_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_10778_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_10788_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_10798_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_10808_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_10818_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_10828_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_10838_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_10848_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_10858_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_10868_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_10878_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_10888_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_10896_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_10904_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_10912_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_10920_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_10928_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_10936_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_10944_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_10952_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_10960_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_10968_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_10976_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_10984_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_10992_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11000_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11008_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11016_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11024_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11032_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11040_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11048_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11056_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11064_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11072_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11080_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11088_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11096_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11104_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11112_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11120_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11128_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11136_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11144_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11152_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11160_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11168_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11176_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11184_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11192_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11200_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11208_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11216_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11224_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11232_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11240_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11248_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11256_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11264_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11272_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11280_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11288_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11296_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11304_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11312_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11320_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11328_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11336_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11344_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11352_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11360_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11368_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11376_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11384_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11392_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11400_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11408_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11416_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11424_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11432_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11440_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11448_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11456_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11464_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11472_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11480_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11488_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11496_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11504_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11512_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11520_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11528_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11536_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11544_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11552_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11560_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11568_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11576_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11584_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11592_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11600_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11608_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11616_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11624_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11632_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11640_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11648_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11656_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11664_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11672_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11680_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11688_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11696_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11704_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11712_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11720_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11728_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11736_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11744_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11752_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11760_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11768_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11776_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11784_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11792_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11800_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11808_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11816_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11824_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11832_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11840_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11848_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11856_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11864_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11872_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11880_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11888_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_11896_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9608_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9618_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9628_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9638_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9648_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9658_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9668_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9678_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9688_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9698_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9708_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9718_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9728_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9738_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9748_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9758_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9768_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9778_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9788_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9798_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9808_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9818_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9828_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9838_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9848_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9858_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9868_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9878_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9888_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9898_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9908_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9918_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9928_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9938_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9948_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9958_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9968_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9978_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9988_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u8_u1_9998_wire : std_logic_vector(0 downto 0);
    signal MA0_9614 : std_logic_vector(7 downto 0);
    signal MA100_10614 : std_logic_vector(7 downto 0);
    signal MA101_10624 : std_logic_vector(7 downto 0);
    signal MA102_10634 : std_logic_vector(7 downto 0);
    signal MA103_10644 : std_logic_vector(7 downto 0);
    signal MA104_10654 : std_logic_vector(7 downto 0);
    signal MA105_10664 : std_logic_vector(7 downto 0);
    signal MA106_10674 : std_logic_vector(7 downto 0);
    signal MA107_10684 : std_logic_vector(7 downto 0);
    signal MA108_10694 : std_logic_vector(7 downto 0);
    signal MA109_10704 : std_logic_vector(7 downto 0);
    signal MA10_9714 : std_logic_vector(7 downto 0);
    signal MA110_10714 : std_logic_vector(7 downto 0);
    signal MA111_10724 : std_logic_vector(7 downto 0);
    signal MA112_10734 : std_logic_vector(7 downto 0);
    signal MA113_10744 : std_logic_vector(7 downto 0);
    signal MA114_10754 : std_logic_vector(7 downto 0);
    signal MA115_10764 : std_logic_vector(7 downto 0);
    signal MA116_10774 : std_logic_vector(7 downto 0);
    signal MA117_10784 : std_logic_vector(7 downto 0);
    signal MA118_10794 : std_logic_vector(7 downto 0);
    signal MA119_10804 : std_logic_vector(7 downto 0);
    signal MA11_9724 : std_logic_vector(7 downto 0);
    signal MA120_10814 : std_logic_vector(7 downto 0);
    signal MA121_10824 : std_logic_vector(7 downto 0);
    signal MA122_10834 : std_logic_vector(7 downto 0);
    signal MA123_10844 : std_logic_vector(7 downto 0);
    signal MA124_10854 : std_logic_vector(7 downto 0);
    signal MA125_10864 : std_logic_vector(7 downto 0);
    signal MA126_10874 : std_logic_vector(7 downto 0);
    signal MA127_10884 : std_logic_vector(7 downto 0);
    signal MA12_9734 : std_logic_vector(7 downto 0);
    signal MA13_9744 : std_logic_vector(7 downto 0);
    signal MA14_9754 : std_logic_vector(7 downto 0);
    signal MA15_9764 : std_logic_vector(7 downto 0);
    signal MA16_9774 : std_logic_vector(7 downto 0);
    signal MA17_9784 : std_logic_vector(7 downto 0);
    signal MA18_9794 : std_logic_vector(7 downto 0);
    signal MA19_9804 : std_logic_vector(7 downto 0);
    signal MA1_9624 : std_logic_vector(7 downto 0);
    signal MA20_9814 : std_logic_vector(7 downto 0);
    signal MA21_9824 : std_logic_vector(7 downto 0);
    signal MA22_9834 : std_logic_vector(7 downto 0);
    signal MA23_9844 : std_logic_vector(7 downto 0);
    signal MA24_9854 : std_logic_vector(7 downto 0);
    signal MA25_9864 : std_logic_vector(7 downto 0);
    signal MA26_9874 : std_logic_vector(7 downto 0);
    signal MA27_9884 : std_logic_vector(7 downto 0);
    signal MA28_9894 : std_logic_vector(7 downto 0);
    signal MA29_9904 : std_logic_vector(7 downto 0);
    signal MA2_9634 : std_logic_vector(7 downto 0);
    signal MA30_9914 : std_logic_vector(7 downto 0);
    signal MA31_9924 : std_logic_vector(7 downto 0);
    signal MA32_9934 : std_logic_vector(7 downto 0);
    signal MA33_9944 : std_logic_vector(7 downto 0);
    signal MA34_9954 : std_logic_vector(7 downto 0);
    signal MA35_9964 : std_logic_vector(7 downto 0);
    signal MA36_9974 : std_logic_vector(7 downto 0);
    signal MA37_9984 : std_logic_vector(7 downto 0);
    signal MA38_9994 : std_logic_vector(7 downto 0);
    signal MA39_10004 : std_logic_vector(7 downto 0);
    signal MA3_9644 : std_logic_vector(7 downto 0);
    signal MA40_10014 : std_logic_vector(7 downto 0);
    signal MA41_10024 : std_logic_vector(7 downto 0);
    signal MA42_10034 : std_logic_vector(7 downto 0);
    signal MA43_10044 : std_logic_vector(7 downto 0);
    signal MA44_10054 : std_logic_vector(7 downto 0);
    signal MA45_10064 : std_logic_vector(7 downto 0);
    signal MA46_10074 : std_logic_vector(7 downto 0);
    signal MA47_10084 : std_logic_vector(7 downto 0);
    signal MA48_10094 : std_logic_vector(7 downto 0);
    signal MA49_10104 : std_logic_vector(7 downto 0);
    signal MA4_9654 : std_logic_vector(7 downto 0);
    signal MA50_10114 : std_logic_vector(7 downto 0);
    signal MA51_10124 : std_logic_vector(7 downto 0);
    signal MA52_10134 : std_logic_vector(7 downto 0);
    signal MA53_10144 : std_logic_vector(7 downto 0);
    signal MA54_10154 : std_logic_vector(7 downto 0);
    signal MA55_10164 : std_logic_vector(7 downto 0);
    signal MA56_10174 : std_logic_vector(7 downto 0);
    signal MA57_10184 : std_logic_vector(7 downto 0);
    signal MA58_10194 : std_logic_vector(7 downto 0);
    signal MA59_10204 : std_logic_vector(7 downto 0);
    signal MA5_9664 : std_logic_vector(7 downto 0);
    signal MA60_10214 : std_logic_vector(7 downto 0);
    signal MA61_10224 : std_logic_vector(7 downto 0);
    signal MA62_10234 : std_logic_vector(7 downto 0);
    signal MA63_10244 : std_logic_vector(7 downto 0);
    signal MA64_10254 : std_logic_vector(7 downto 0);
    signal MA65_10264 : std_logic_vector(7 downto 0);
    signal MA66_10274 : std_logic_vector(7 downto 0);
    signal MA67_10284 : std_logic_vector(7 downto 0);
    signal MA68_10294 : std_logic_vector(7 downto 0);
    signal MA69_10304 : std_logic_vector(7 downto 0);
    signal MA6_9674 : std_logic_vector(7 downto 0);
    signal MA70_10314 : std_logic_vector(7 downto 0);
    signal MA71_10324 : std_logic_vector(7 downto 0);
    signal MA72_10334 : std_logic_vector(7 downto 0);
    signal MA73_10344 : std_logic_vector(7 downto 0);
    signal MA74_10354 : std_logic_vector(7 downto 0);
    signal MA75_10364 : std_logic_vector(7 downto 0);
    signal MA76_10374 : std_logic_vector(7 downto 0);
    signal MA77_10384 : std_logic_vector(7 downto 0);
    signal MA78_10394 : std_logic_vector(7 downto 0);
    signal MA79_10404 : std_logic_vector(7 downto 0);
    signal MA7_9684 : std_logic_vector(7 downto 0);
    signal MA80_10414 : std_logic_vector(7 downto 0);
    signal MA81_10424 : std_logic_vector(7 downto 0);
    signal MA82_10434 : std_logic_vector(7 downto 0);
    signal MA83_10444 : std_logic_vector(7 downto 0);
    signal MA84_10454 : std_logic_vector(7 downto 0);
    signal MA85_10464 : std_logic_vector(7 downto 0);
    signal MA86_10474 : std_logic_vector(7 downto 0);
    signal MA87_10484 : std_logic_vector(7 downto 0);
    signal MA88_10494 : std_logic_vector(7 downto 0);
    signal MA89_10504 : std_logic_vector(7 downto 0);
    signal MA8_9694 : std_logic_vector(7 downto 0);
    signal MA90_10514 : std_logic_vector(7 downto 0);
    signal MA91_10524 : std_logic_vector(7 downto 0);
    signal MA92_10534 : std_logic_vector(7 downto 0);
    signal MA93_10544 : std_logic_vector(7 downto 0);
    signal MA94_10554 : std_logic_vector(7 downto 0);
    signal MA95_10564 : std_logic_vector(7 downto 0);
    signal MA96_10574 : std_logic_vector(7 downto 0);
    signal MA97_10584 : std_logic_vector(7 downto 0);
    signal MA98_10594 : std_logic_vector(7 downto 0);
    signal MA99_10604 : std_logic_vector(7 downto 0);
    signal MA9_9704 : std_logic_vector(7 downto 0);
    signal MB0_10892 : std_logic_vector(7 downto 0);
    signal MB10_10972 : std_logic_vector(7 downto 0);
    signal MB11_10980 : std_logic_vector(7 downto 0);
    signal MB12_10988 : std_logic_vector(7 downto 0);
    signal MB13_10996 : std_logic_vector(7 downto 0);
    signal MB14_11004 : std_logic_vector(7 downto 0);
    signal MB15_11012 : std_logic_vector(7 downto 0);
    signal MB16_11020 : std_logic_vector(7 downto 0);
    signal MB17_11028 : std_logic_vector(7 downto 0);
    signal MB18_11036 : std_logic_vector(7 downto 0);
    signal MB19_11044 : std_logic_vector(7 downto 0);
    signal MB1_10900 : std_logic_vector(7 downto 0);
    signal MB20_11052 : std_logic_vector(7 downto 0);
    signal MB21_11060 : std_logic_vector(7 downto 0);
    signal MB22_11068 : std_logic_vector(7 downto 0);
    signal MB23_11076 : std_logic_vector(7 downto 0);
    signal MB24_11084 : std_logic_vector(7 downto 0);
    signal MB25_11092 : std_logic_vector(7 downto 0);
    signal MB26_11100 : std_logic_vector(7 downto 0);
    signal MB27_11108 : std_logic_vector(7 downto 0);
    signal MB28_11116 : std_logic_vector(7 downto 0);
    signal MB29_11124 : std_logic_vector(7 downto 0);
    signal MB2_10908 : std_logic_vector(7 downto 0);
    signal MB30_11132 : std_logic_vector(7 downto 0);
    signal MB31_11140 : std_logic_vector(7 downto 0);
    signal MB32_11148 : std_logic_vector(7 downto 0);
    signal MB33_11156 : std_logic_vector(7 downto 0);
    signal MB34_11164 : std_logic_vector(7 downto 0);
    signal MB35_11172 : std_logic_vector(7 downto 0);
    signal MB36_11180 : std_logic_vector(7 downto 0);
    signal MB37_11188 : std_logic_vector(7 downto 0);
    signal MB38_11196 : std_logic_vector(7 downto 0);
    signal MB39_11204 : std_logic_vector(7 downto 0);
    signal MB3_10916 : std_logic_vector(7 downto 0);
    signal MB40_11212 : std_logic_vector(7 downto 0);
    signal MB41_11220 : std_logic_vector(7 downto 0);
    signal MB42_11228 : std_logic_vector(7 downto 0);
    signal MB43_11236 : std_logic_vector(7 downto 0);
    signal MB44_11244 : std_logic_vector(7 downto 0);
    signal MB45_11252 : std_logic_vector(7 downto 0);
    signal MB46_11260 : std_logic_vector(7 downto 0);
    signal MB47_11268 : std_logic_vector(7 downto 0);
    signal MB48_11276 : std_logic_vector(7 downto 0);
    signal MB49_11284 : std_logic_vector(7 downto 0);
    signal MB4_10924 : std_logic_vector(7 downto 0);
    signal MB50_11292 : std_logic_vector(7 downto 0);
    signal MB51_11300 : std_logic_vector(7 downto 0);
    signal MB52_11308 : std_logic_vector(7 downto 0);
    signal MB53_11316 : std_logic_vector(7 downto 0);
    signal MB54_11324 : std_logic_vector(7 downto 0);
    signal MB55_11332 : std_logic_vector(7 downto 0);
    signal MB56_11340 : std_logic_vector(7 downto 0);
    signal MB57_11348 : std_logic_vector(7 downto 0);
    signal MB58_11356 : std_logic_vector(7 downto 0);
    signal MB59_11364 : std_logic_vector(7 downto 0);
    signal MB5_10932 : std_logic_vector(7 downto 0);
    signal MB60_11372 : std_logic_vector(7 downto 0);
    signal MB61_11380 : std_logic_vector(7 downto 0);
    signal MB62_11388 : std_logic_vector(7 downto 0);
    signal MB63_11396 : std_logic_vector(7 downto 0);
    signal MB6_10940 : std_logic_vector(7 downto 0);
    signal MB7_10948 : std_logic_vector(7 downto 0);
    signal MB8_10956 : std_logic_vector(7 downto 0);
    signal MB9_10964 : std_logic_vector(7 downto 0);
    signal MC0_11404 : std_logic_vector(7 downto 0);
    signal MC10_11484 : std_logic_vector(7 downto 0);
    signal MC11_11492 : std_logic_vector(7 downto 0);
    signal MC12_11500 : std_logic_vector(7 downto 0);
    signal MC13_11508 : std_logic_vector(7 downto 0);
    signal MC14_11516 : std_logic_vector(7 downto 0);
    signal MC15_11524 : std_logic_vector(7 downto 0);
    signal MC16_11532 : std_logic_vector(7 downto 0);
    signal MC17_11540 : std_logic_vector(7 downto 0);
    signal MC18_11548 : std_logic_vector(7 downto 0);
    signal MC19_11556 : std_logic_vector(7 downto 0);
    signal MC1_11412 : std_logic_vector(7 downto 0);
    signal MC20_11564 : std_logic_vector(7 downto 0);
    signal MC21_11572 : std_logic_vector(7 downto 0);
    signal MC22_11580 : std_logic_vector(7 downto 0);
    signal MC23_11588 : std_logic_vector(7 downto 0);
    signal MC24_11596 : std_logic_vector(7 downto 0);
    signal MC25_11604 : std_logic_vector(7 downto 0);
    signal MC26_11612 : std_logic_vector(7 downto 0);
    signal MC27_11620 : std_logic_vector(7 downto 0);
    signal MC28_11628 : std_logic_vector(7 downto 0);
    signal MC29_11636 : std_logic_vector(7 downto 0);
    signal MC2_11420 : std_logic_vector(7 downto 0);
    signal MC30_11644 : std_logic_vector(7 downto 0);
    signal MC31_11652 : std_logic_vector(7 downto 0);
    signal MC3_11428 : std_logic_vector(7 downto 0);
    signal MC4_11436 : std_logic_vector(7 downto 0);
    signal MC5_11444 : std_logic_vector(7 downto 0);
    signal MC6_11452 : std_logic_vector(7 downto 0);
    signal MC7_11460 : std_logic_vector(7 downto 0);
    signal MC8_11468 : std_logic_vector(7 downto 0);
    signal MC9_11476 : std_logic_vector(7 downto 0);
    signal MD0_11660 : std_logic_vector(7 downto 0);
    signal MD10_11740 : std_logic_vector(7 downto 0);
    signal MD11_11748 : std_logic_vector(7 downto 0);
    signal MD12_11756 : std_logic_vector(7 downto 0);
    signal MD13_11764 : std_logic_vector(7 downto 0);
    signal MD14_11772 : std_logic_vector(7 downto 0);
    signal MD15_11780 : std_logic_vector(7 downto 0);
    signal MD1_11668 : std_logic_vector(7 downto 0);
    signal MD2_11676 : std_logic_vector(7 downto 0);
    signal MD3_11684 : std_logic_vector(7 downto 0);
    signal MD4_11692 : std_logic_vector(7 downto 0);
    signal MD5_11700 : std_logic_vector(7 downto 0);
    signal MD6_11708 : std_logic_vector(7 downto 0);
    signal MD7_11716 : std_logic_vector(7 downto 0);
    signal MD8_11724 : std_logic_vector(7 downto 0);
    signal MD9_11732 : std_logic_vector(7 downto 0);
    signal ME0_11788 : std_logic_vector(7 downto 0);
    signal ME1_11796 : std_logic_vector(7 downto 0);
    signal ME2_11804 : std_logic_vector(7 downto 0);
    signal ME3_11812 : std_logic_vector(7 downto 0);
    signal ME4_11820 : std_logic_vector(7 downto 0);
    signal ME5_11828 : std_logic_vector(7 downto 0);
    signal ME6_11836 : std_logic_vector(7 downto 0);
    signal ME7_11844 : std_logic_vector(7 downto 0);
    signal MF0_11852 : std_logic_vector(7 downto 0);
    signal MF1_11860 : std_logic_vector(7 downto 0);
    signal MF2_11868 : std_logic_vector(7 downto 0);
    signal MF3_11876 : std_logic_vector(7 downto 0);
    signal MG0_11884 : std_logic_vector(7 downto 0);
    signal MG1_11892 : std_logic_vector(7 downto 0);
    signal konst_10007_wire_constant : std_logic_vector(7 downto 0);
    signal konst_10017_wire_constant : std_logic_vector(7 downto 0);
    signal konst_10027_wire_constant : std_logic_vector(7 downto 0);
    signal konst_10037_wire_constant : std_logic_vector(7 downto 0);
    signal konst_10047_wire_constant : std_logic_vector(7 downto 0);
    signal konst_10057_wire_constant : std_logic_vector(7 downto 0);
    signal konst_10067_wire_constant : std_logic_vector(7 downto 0);
    signal konst_10077_wire_constant : std_logic_vector(7 downto 0);
    signal konst_10087_wire_constant : std_logic_vector(7 downto 0);
    signal konst_10097_wire_constant : std_logic_vector(7 downto 0);
    signal konst_10107_wire_constant : std_logic_vector(7 downto 0);
    signal konst_10117_wire_constant : std_logic_vector(7 downto 0);
    signal konst_10127_wire_constant : std_logic_vector(7 downto 0);
    signal konst_10137_wire_constant : std_logic_vector(7 downto 0);
    signal konst_10147_wire_constant : std_logic_vector(7 downto 0);
    signal konst_10157_wire_constant : std_logic_vector(7 downto 0);
    signal konst_10167_wire_constant : std_logic_vector(7 downto 0);
    signal konst_10177_wire_constant : std_logic_vector(7 downto 0);
    signal konst_10187_wire_constant : std_logic_vector(7 downto 0);
    signal konst_10197_wire_constant : std_logic_vector(7 downto 0);
    signal konst_10207_wire_constant : std_logic_vector(7 downto 0);
    signal konst_10217_wire_constant : std_logic_vector(7 downto 0);
    signal konst_10227_wire_constant : std_logic_vector(7 downto 0);
    signal konst_10237_wire_constant : std_logic_vector(7 downto 0);
    signal konst_10247_wire_constant : std_logic_vector(7 downto 0);
    signal konst_10257_wire_constant : std_logic_vector(7 downto 0);
    signal konst_10267_wire_constant : std_logic_vector(7 downto 0);
    signal konst_10277_wire_constant : std_logic_vector(7 downto 0);
    signal konst_10287_wire_constant : std_logic_vector(7 downto 0);
    signal konst_10297_wire_constant : std_logic_vector(7 downto 0);
    signal konst_10307_wire_constant : std_logic_vector(7 downto 0);
    signal konst_10317_wire_constant : std_logic_vector(7 downto 0);
    signal konst_10327_wire_constant : std_logic_vector(7 downto 0);
    signal konst_10337_wire_constant : std_logic_vector(7 downto 0);
    signal konst_10347_wire_constant : std_logic_vector(7 downto 0);
    signal konst_10357_wire_constant : std_logic_vector(7 downto 0);
    signal konst_10367_wire_constant : std_logic_vector(7 downto 0);
    signal konst_10377_wire_constant : std_logic_vector(7 downto 0);
    signal konst_10387_wire_constant : std_logic_vector(7 downto 0);
    signal konst_10397_wire_constant : std_logic_vector(7 downto 0);
    signal konst_10407_wire_constant : std_logic_vector(7 downto 0);
    signal konst_10417_wire_constant : std_logic_vector(7 downto 0);
    signal konst_10427_wire_constant : std_logic_vector(7 downto 0);
    signal konst_10437_wire_constant : std_logic_vector(7 downto 0);
    signal konst_10447_wire_constant : std_logic_vector(7 downto 0);
    signal konst_10457_wire_constant : std_logic_vector(7 downto 0);
    signal konst_10467_wire_constant : std_logic_vector(7 downto 0);
    signal konst_10477_wire_constant : std_logic_vector(7 downto 0);
    signal konst_10487_wire_constant : std_logic_vector(7 downto 0);
    signal konst_10497_wire_constant : std_logic_vector(7 downto 0);
    signal konst_10507_wire_constant : std_logic_vector(7 downto 0);
    signal konst_10517_wire_constant : std_logic_vector(7 downto 0);
    signal konst_10527_wire_constant : std_logic_vector(7 downto 0);
    signal konst_10537_wire_constant : std_logic_vector(7 downto 0);
    signal konst_10547_wire_constant : std_logic_vector(7 downto 0);
    signal konst_10557_wire_constant : std_logic_vector(7 downto 0);
    signal konst_10567_wire_constant : std_logic_vector(7 downto 0);
    signal konst_10577_wire_constant : std_logic_vector(7 downto 0);
    signal konst_10587_wire_constant : std_logic_vector(7 downto 0);
    signal konst_10597_wire_constant : std_logic_vector(7 downto 0);
    signal konst_10607_wire_constant : std_logic_vector(7 downto 0);
    signal konst_10617_wire_constant : std_logic_vector(7 downto 0);
    signal konst_10627_wire_constant : std_logic_vector(7 downto 0);
    signal konst_10637_wire_constant : std_logic_vector(7 downto 0);
    signal konst_10647_wire_constant : std_logic_vector(7 downto 0);
    signal konst_10657_wire_constant : std_logic_vector(7 downto 0);
    signal konst_10667_wire_constant : std_logic_vector(7 downto 0);
    signal konst_10677_wire_constant : std_logic_vector(7 downto 0);
    signal konst_10687_wire_constant : std_logic_vector(7 downto 0);
    signal konst_10697_wire_constant : std_logic_vector(7 downto 0);
    signal konst_10707_wire_constant : std_logic_vector(7 downto 0);
    signal konst_10717_wire_constant : std_logic_vector(7 downto 0);
    signal konst_10727_wire_constant : std_logic_vector(7 downto 0);
    signal konst_10737_wire_constant : std_logic_vector(7 downto 0);
    signal konst_10747_wire_constant : std_logic_vector(7 downto 0);
    signal konst_10757_wire_constant : std_logic_vector(7 downto 0);
    signal konst_10767_wire_constant : std_logic_vector(7 downto 0);
    signal konst_10777_wire_constant : std_logic_vector(7 downto 0);
    signal konst_10787_wire_constant : std_logic_vector(7 downto 0);
    signal konst_10797_wire_constant : std_logic_vector(7 downto 0);
    signal konst_10807_wire_constant : std_logic_vector(7 downto 0);
    signal konst_10817_wire_constant : std_logic_vector(7 downto 0);
    signal konst_10827_wire_constant : std_logic_vector(7 downto 0);
    signal konst_10837_wire_constant : std_logic_vector(7 downto 0);
    signal konst_10847_wire_constant : std_logic_vector(7 downto 0);
    signal konst_10857_wire_constant : std_logic_vector(7 downto 0);
    signal konst_10867_wire_constant : std_logic_vector(7 downto 0);
    signal konst_10877_wire_constant : std_logic_vector(7 downto 0);
    signal konst_10887_wire_constant : std_logic_vector(7 downto 0);
    signal konst_10895_wire_constant : std_logic_vector(7 downto 0);
    signal konst_10903_wire_constant : std_logic_vector(7 downto 0);
    signal konst_10911_wire_constant : std_logic_vector(7 downto 0);
    signal konst_10919_wire_constant : std_logic_vector(7 downto 0);
    signal konst_10927_wire_constant : std_logic_vector(7 downto 0);
    signal konst_10935_wire_constant : std_logic_vector(7 downto 0);
    signal konst_10943_wire_constant : std_logic_vector(7 downto 0);
    signal konst_10951_wire_constant : std_logic_vector(7 downto 0);
    signal konst_10959_wire_constant : std_logic_vector(7 downto 0);
    signal konst_10967_wire_constant : std_logic_vector(7 downto 0);
    signal konst_10975_wire_constant : std_logic_vector(7 downto 0);
    signal konst_10983_wire_constant : std_logic_vector(7 downto 0);
    signal konst_10991_wire_constant : std_logic_vector(7 downto 0);
    signal konst_10999_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11007_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11015_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11023_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11031_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11039_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11047_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11055_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11063_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11071_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11079_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11087_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11095_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11103_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11111_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11119_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11127_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11135_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11143_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11151_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11159_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11167_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11175_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11183_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11191_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11199_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11207_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11215_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11223_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11231_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11239_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11247_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11255_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11263_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11271_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11279_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11287_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11295_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11303_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11311_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11319_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11327_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11335_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11343_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11351_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11359_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11367_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11375_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11383_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11391_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11399_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11407_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11415_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11423_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11431_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11439_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11447_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11455_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11463_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11471_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11479_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11487_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11495_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11503_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11511_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11519_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11527_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11535_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11543_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11551_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11559_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11567_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11575_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11583_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11591_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11599_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11607_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11615_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11623_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11631_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11639_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11647_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11655_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11663_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11671_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11679_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11687_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11695_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11703_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11711_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11719_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11727_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11735_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11743_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11751_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11759_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11767_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11775_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11783_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11791_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11799_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11807_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11815_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11823_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11831_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11839_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11847_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11855_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11863_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11871_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11879_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11887_wire_constant : std_logic_vector(7 downto 0);
    signal konst_11895_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9607_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9617_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9627_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9637_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9647_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9657_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9667_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9677_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9687_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9697_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9707_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9717_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9727_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9737_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9747_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9757_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9767_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9777_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9787_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9797_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9807_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9817_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9827_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9837_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9847_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9857_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9867_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9877_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9887_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9897_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9907_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9917_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9927_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9937_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9947_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9957_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9967_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9977_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9987_wire_constant : std_logic_vector(7 downto 0);
    signal konst_9997_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10000_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10002_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10010_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10012_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10020_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10022_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10030_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10032_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10040_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10042_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10050_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10052_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10060_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10062_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10070_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10072_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10080_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10082_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10090_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10092_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10100_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10102_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10110_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10112_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10120_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10122_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10130_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10132_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10140_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10142_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10150_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10152_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10160_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10162_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10170_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10172_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10180_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10182_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10190_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10192_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10200_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10202_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10210_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10212_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10220_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10222_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10230_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10232_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10240_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10242_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10250_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10252_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10260_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10262_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10270_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10272_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10280_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10282_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10290_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10292_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10300_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10302_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10310_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10312_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10320_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10322_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10330_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10332_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10340_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10342_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10350_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10352_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10360_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10362_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10370_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10372_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10380_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10382_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10390_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10392_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10400_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10402_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10410_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10412_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10420_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10422_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10430_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10432_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10440_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10442_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10450_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10452_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10460_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10462_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10470_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10472_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10480_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10482_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10490_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10492_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10500_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10502_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10510_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10512_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10520_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10522_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10530_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10532_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10540_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10542_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10550_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10552_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10560_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10562_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10570_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10572_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10580_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10582_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10590_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10592_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10600_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10602_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10610_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10612_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10620_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10622_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10630_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10632_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10640_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10642_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10650_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10652_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10660_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10662_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10670_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10672_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10680_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10682_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10690_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10692_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10700_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10702_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10710_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10712_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10720_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10722_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10730_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10732_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10740_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10742_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10750_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10752_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10760_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10762_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10770_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10772_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10780_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10782_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10790_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10792_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10800_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10802_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10810_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10812_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10820_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10822_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10830_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10832_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10840_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10842_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10850_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10852_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10860_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10862_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10870_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10872_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10880_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_10882_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_9610_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_9612_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_9620_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_9622_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_9630_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_9632_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_9640_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_9642_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_9650_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_9652_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_9660_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_9662_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_9670_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_9672_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_9680_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_9682_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_9690_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_9692_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_9700_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_9702_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_9710_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_9712_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_9720_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_9722_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_9730_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_9732_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_9740_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_9742_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_9750_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_9752_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_9760_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_9762_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_9770_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_9772_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_9780_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_9782_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_9790_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_9792_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_9800_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_9802_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_9810_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_9812_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_9820_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_9822_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_9830_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_9832_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_9840_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_9842_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_9850_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_9852_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_9860_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_9862_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_9870_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_9872_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_9880_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_9882_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_9890_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_9892_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_9900_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_9902_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_9910_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_9912_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_9920_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_9922_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_9930_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_9932_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_9940_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_9942_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_9950_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_9952_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_9960_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_9962_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_9970_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_9972_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_9980_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_9982_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_9990_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_9992_wire_constant : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    konst_10007_wire_constant <= "00000000";
    konst_10017_wire_constant <= "00000000";
    konst_10027_wire_constant <= "00000000";
    konst_10037_wire_constant <= "00000000";
    konst_10047_wire_constant <= "00000000";
    konst_10057_wire_constant <= "00000000";
    konst_10067_wire_constant <= "00000000";
    konst_10077_wire_constant <= "00000000";
    konst_10087_wire_constant <= "00000000";
    konst_10097_wire_constant <= "00000000";
    konst_10107_wire_constant <= "00000000";
    konst_10117_wire_constant <= "00000000";
    konst_10127_wire_constant <= "00000000";
    konst_10137_wire_constant <= "00000000";
    konst_10147_wire_constant <= "00000000";
    konst_10157_wire_constant <= "00000000";
    konst_10167_wire_constant <= "00000000";
    konst_10177_wire_constant <= "00000000";
    konst_10187_wire_constant <= "00000000";
    konst_10197_wire_constant <= "00000000";
    konst_10207_wire_constant <= "00000000";
    konst_10217_wire_constant <= "00000000";
    konst_10227_wire_constant <= "00000000";
    konst_10237_wire_constant <= "00000000";
    konst_10247_wire_constant <= "00000000";
    konst_10257_wire_constant <= "00000000";
    konst_10267_wire_constant <= "00000000";
    konst_10277_wire_constant <= "00000000";
    konst_10287_wire_constant <= "00000000";
    konst_10297_wire_constant <= "00000000";
    konst_10307_wire_constant <= "00000000";
    konst_10317_wire_constant <= "00000000";
    konst_10327_wire_constant <= "00000000";
    konst_10337_wire_constant <= "00000000";
    konst_10347_wire_constant <= "00000000";
    konst_10357_wire_constant <= "00000000";
    konst_10367_wire_constant <= "00000000";
    konst_10377_wire_constant <= "00000000";
    konst_10387_wire_constant <= "00000000";
    konst_10397_wire_constant <= "00000000";
    konst_10407_wire_constant <= "00000000";
    konst_10417_wire_constant <= "00000000";
    konst_10427_wire_constant <= "00000000";
    konst_10437_wire_constant <= "00000000";
    konst_10447_wire_constant <= "00000000";
    konst_10457_wire_constant <= "00000000";
    konst_10467_wire_constant <= "00000000";
    konst_10477_wire_constant <= "00000000";
    konst_10487_wire_constant <= "00000000";
    konst_10497_wire_constant <= "00000000";
    konst_10507_wire_constant <= "00000000";
    konst_10517_wire_constant <= "00000000";
    konst_10527_wire_constant <= "00000000";
    konst_10537_wire_constant <= "00000000";
    konst_10547_wire_constant <= "00000000";
    konst_10557_wire_constant <= "00000000";
    konst_10567_wire_constant <= "00000000";
    konst_10577_wire_constant <= "00000000";
    konst_10587_wire_constant <= "00000000";
    konst_10597_wire_constant <= "00000000";
    konst_10607_wire_constant <= "00000000";
    konst_10617_wire_constant <= "00000000";
    konst_10627_wire_constant <= "00000000";
    konst_10637_wire_constant <= "00000000";
    konst_10647_wire_constant <= "00000000";
    konst_10657_wire_constant <= "00000000";
    konst_10667_wire_constant <= "00000000";
    konst_10677_wire_constant <= "00000000";
    konst_10687_wire_constant <= "00000000";
    konst_10697_wire_constant <= "00000000";
    konst_10707_wire_constant <= "00000000";
    konst_10717_wire_constant <= "00000000";
    konst_10727_wire_constant <= "00000000";
    konst_10737_wire_constant <= "00000000";
    konst_10747_wire_constant <= "00000000";
    konst_10757_wire_constant <= "00000000";
    konst_10767_wire_constant <= "00000000";
    konst_10777_wire_constant <= "00000000";
    konst_10787_wire_constant <= "00000000";
    konst_10797_wire_constant <= "00000000";
    konst_10807_wire_constant <= "00000000";
    konst_10817_wire_constant <= "00000000";
    konst_10827_wire_constant <= "00000000";
    konst_10837_wire_constant <= "00000000";
    konst_10847_wire_constant <= "00000000";
    konst_10857_wire_constant <= "00000000";
    konst_10867_wire_constant <= "00000000";
    konst_10877_wire_constant <= "00000000";
    konst_10887_wire_constant <= "00000001";
    konst_10895_wire_constant <= "00000001";
    konst_10903_wire_constant <= "00000001";
    konst_10911_wire_constant <= "00000001";
    konst_10919_wire_constant <= "00000001";
    konst_10927_wire_constant <= "00000001";
    konst_10935_wire_constant <= "00000001";
    konst_10943_wire_constant <= "00000001";
    konst_10951_wire_constant <= "00000001";
    konst_10959_wire_constant <= "00000001";
    konst_10967_wire_constant <= "00000001";
    konst_10975_wire_constant <= "00000001";
    konst_10983_wire_constant <= "00000001";
    konst_10991_wire_constant <= "00000001";
    konst_10999_wire_constant <= "00000001";
    konst_11007_wire_constant <= "00000001";
    konst_11015_wire_constant <= "00000001";
    konst_11023_wire_constant <= "00000001";
    konst_11031_wire_constant <= "00000001";
    konst_11039_wire_constant <= "00000001";
    konst_11047_wire_constant <= "00000001";
    konst_11055_wire_constant <= "00000001";
    konst_11063_wire_constant <= "00000001";
    konst_11071_wire_constant <= "00000001";
    konst_11079_wire_constant <= "00000001";
    konst_11087_wire_constant <= "00000001";
    konst_11095_wire_constant <= "00000001";
    konst_11103_wire_constant <= "00000001";
    konst_11111_wire_constant <= "00000001";
    konst_11119_wire_constant <= "00000001";
    konst_11127_wire_constant <= "00000001";
    konst_11135_wire_constant <= "00000001";
    konst_11143_wire_constant <= "00000001";
    konst_11151_wire_constant <= "00000001";
    konst_11159_wire_constant <= "00000001";
    konst_11167_wire_constant <= "00000001";
    konst_11175_wire_constant <= "00000001";
    konst_11183_wire_constant <= "00000001";
    konst_11191_wire_constant <= "00000001";
    konst_11199_wire_constant <= "00000001";
    konst_11207_wire_constant <= "00000001";
    konst_11215_wire_constant <= "00000001";
    konst_11223_wire_constant <= "00000001";
    konst_11231_wire_constant <= "00000001";
    konst_11239_wire_constant <= "00000001";
    konst_11247_wire_constant <= "00000001";
    konst_11255_wire_constant <= "00000001";
    konst_11263_wire_constant <= "00000001";
    konst_11271_wire_constant <= "00000001";
    konst_11279_wire_constant <= "00000001";
    konst_11287_wire_constant <= "00000001";
    konst_11295_wire_constant <= "00000001";
    konst_11303_wire_constant <= "00000001";
    konst_11311_wire_constant <= "00000001";
    konst_11319_wire_constant <= "00000001";
    konst_11327_wire_constant <= "00000001";
    konst_11335_wire_constant <= "00000001";
    konst_11343_wire_constant <= "00000001";
    konst_11351_wire_constant <= "00000001";
    konst_11359_wire_constant <= "00000001";
    konst_11367_wire_constant <= "00000001";
    konst_11375_wire_constant <= "00000001";
    konst_11383_wire_constant <= "00000001";
    konst_11391_wire_constant <= "00000001";
    konst_11399_wire_constant <= "00000010";
    konst_11407_wire_constant <= "00000010";
    konst_11415_wire_constant <= "00000010";
    konst_11423_wire_constant <= "00000010";
    konst_11431_wire_constant <= "00000010";
    konst_11439_wire_constant <= "00000010";
    konst_11447_wire_constant <= "00000010";
    konst_11455_wire_constant <= "00000010";
    konst_11463_wire_constant <= "00000010";
    konst_11471_wire_constant <= "00000010";
    konst_11479_wire_constant <= "00000010";
    konst_11487_wire_constant <= "00000010";
    konst_11495_wire_constant <= "00000010";
    konst_11503_wire_constant <= "00000010";
    konst_11511_wire_constant <= "00000010";
    konst_11519_wire_constant <= "00000010";
    konst_11527_wire_constant <= "00000010";
    konst_11535_wire_constant <= "00000010";
    konst_11543_wire_constant <= "00000010";
    konst_11551_wire_constant <= "00000010";
    konst_11559_wire_constant <= "00000010";
    konst_11567_wire_constant <= "00000010";
    konst_11575_wire_constant <= "00000010";
    konst_11583_wire_constant <= "00000010";
    konst_11591_wire_constant <= "00000010";
    konst_11599_wire_constant <= "00000010";
    konst_11607_wire_constant <= "00000010";
    konst_11615_wire_constant <= "00000010";
    konst_11623_wire_constant <= "00000010";
    konst_11631_wire_constant <= "00000010";
    konst_11639_wire_constant <= "00000010";
    konst_11647_wire_constant <= "00000010";
    konst_11655_wire_constant <= "00000011";
    konst_11663_wire_constant <= "00000011";
    konst_11671_wire_constant <= "00000011";
    konst_11679_wire_constant <= "00000011";
    konst_11687_wire_constant <= "00000011";
    konst_11695_wire_constant <= "00000011";
    konst_11703_wire_constant <= "00000011";
    konst_11711_wire_constant <= "00000011";
    konst_11719_wire_constant <= "00000011";
    konst_11727_wire_constant <= "00000011";
    konst_11735_wire_constant <= "00000011";
    konst_11743_wire_constant <= "00000011";
    konst_11751_wire_constant <= "00000011";
    konst_11759_wire_constant <= "00000011";
    konst_11767_wire_constant <= "00000011";
    konst_11775_wire_constant <= "00000011";
    konst_11783_wire_constant <= "00000100";
    konst_11791_wire_constant <= "00000100";
    konst_11799_wire_constant <= "00000100";
    konst_11807_wire_constant <= "00000100";
    konst_11815_wire_constant <= "00000100";
    konst_11823_wire_constant <= "00000100";
    konst_11831_wire_constant <= "00000100";
    konst_11839_wire_constant <= "00000100";
    konst_11847_wire_constant <= "00000101";
    konst_11855_wire_constant <= "00000101";
    konst_11863_wire_constant <= "00000101";
    konst_11871_wire_constant <= "00000101";
    konst_11879_wire_constant <= "00000110";
    konst_11887_wire_constant <= "00000110";
    konst_11895_wire_constant <= "00000111";
    konst_9607_wire_constant <= "00000000";
    konst_9617_wire_constant <= "00000000";
    konst_9627_wire_constant <= "00000000";
    konst_9637_wire_constant <= "00000000";
    konst_9647_wire_constant <= "00000000";
    konst_9657_wire_constant <= "00000000";
    konst_9667_wire_constant <= "00000000";
    konst_9677_wire_constant <= "00000000";
    konst_9687_wire_constant <= "00000000";
    konst_9697_wire_constant <= "00000000";
    konst_9707_wire_constant <= "00000000";
    konst_9717_wire_constant <= "00000000";
    konst_9727_wire_constant <= "00000000";
    konst_9737_wire_constant <= "00000000";
    konst_9747_wire_constant <= "00000000";
    konst_9757_wire_constant <= "00000000";
    konst_9767_wire_constant <= "00000000";
    konst_9777_wire_constant <= "00000000";
    konst_9787_wire_constant <= "00000000";
    konst_9797_wire_constant <= "00000000";
    konst_9807_wire_constant <= "00000000";
    konst_9817_wire_constant <= "00000000";
    konst_9827_wire_constant <= "00000000";
    konst_9837_wire_constant <= "00000000";
    konst_9847_wire_constant <= "00000000";
    konst_9857_wire_constant <= "00000000";
    konst_9867_wire_constant <= "00000000";
    konst_9877_wire_constant <= "00000000";
    konst_9887_wire_constant <= "00000000";
    konst_9897_wire_constant <= "00000000";
    konst_9907_wire_constant <= "00000000";
    konst_9917_wire_constant <= "00000000";
    konst_9927_wire_constant <= "00000000";
    konst_9937_wire_constant <= "00000000";
    konst_9947_wire_constant <= "00000000";
    konst_9957_wire_constant <= "00000000";
    konst_9967_wire_constant <= "00000000";
    konst_9977_wire_constant <= "00000000";
    konst_9987_wire_constant <= "00000000";
    konst_9997_wire_constant <= "00000000";
    type_cast_10000_wire_constant <= "10000100";
    type_cast_10002_wire_constant <= "00101111";
    type_cast_10010_wire_constant <= "11010001";
    type_cast_10012_wire_constant <= "01010011";
    type_cast_10020_wire_constant <= "11101101";
    type_cast_10022_wire_constant <= "00000000";
    type_cast_10030_wire_constant <= "11111100";
    type_cast_10032_wire_constant <= "00100000";
    type_cast_10040_wire_constant <= "01011011";
    type_cast_10042_wire_constant <= "10110001";
    type_cast_10050_wire_constant <= "11001011";
    type_cast_10052_wire_constant <= "01101010";
    type_cast_10060_wire_constant <= "00111001";
    type_cast_10062_wire_constant <= "10111110";
    type_cast_10070_wire_constant <= "01001100";
    type_cast_10072_wire_constant <= "01001010";
    type_cast_10080_wire_constant <= "11001111";
    type_cast_10082_wire_constant <= "01011000";
    type_cast_10090_wire_constant <= "11101111";
    type_cast_10092_wire_constant <= "11010000";
    type_cast_10100_wire_constant <= "11111011";
    type_cast_10102_wire_constant <= "10101010";
    type_cast_10110_wire_constant <= "01001101";
    type_cast_10112_wire_constant <= "01000011";
    type_cast_10120_wire_constant <= "10000101";
    type_cast_10122_wire_constant <= "00110011";
    type_cast_10130_wire_constant <= "11111001";
    type_cast_10132_wire_constant <= "01000101";
    type_cast_10140_wire_constant <= "01111111";
    type_cast_10142_wire_constant <= "00000010";
    type_cast_10150_wire_constant <= "00111100";
    type_cast_10152_wire_constant <= "01010000";
    type_cast_10160_wire_constant <= "10101000";
    type_cast_10162_wire_constant <= "10011111";
    type_cast_10170_wire_constant <= "10100011";
    type_cast_10172_wire_constant <= "01010001";
    type_cast_10180_wire_constant <= "10001111";
    type_cast_10182_wire_constant <= "01000000";
    type_cast_10190_wire_constant <= "10011101";
    type_cast_10192_wire_constant <= "10010010";
    type_cast_10200_wire_constant <= "11110101";
    type_cast_10202_wire_constant <= "00111000";
    type_cast_10210_wire_constant <= "10110110";
    type_cast_10212_wire_constant <= "10111100";
    type_cast_10220_wire_constant <= "00100001";
    type_cast_10222_wire_constant <= "11011010";
    type_cast_10230_wire_constant <= "11111111";
    type_cast_10232_wire_constant <= "00010000";
    type_cast_10240_wire_constant <= "11010010";
    type_cast_10242_wire_constant <= "11110011";
    type_cast_10250_wire_constant <= "00001100";
    type_cast_10252_wire_constant <= "11001101";
    type_cast_10260_wire_constant <= "11101100";
    type_cast_10262_wire_constant <= "00010011";
    type_cast_10270_wire_constant <= "10010111";
    type_cast_10272_wire_constant <= "01011111";
    type_cast_10280_wire_constant <= "00010111";
    type_cast_10282_wire_constant <= "01000100";
    type_cast_10290_wire_constant <= "10100111";
    type_cast_10292_wire_constant <= "11000100";
    type_cast_10300_wire_constant <= "00111101";
    type_cast_10302_wire_constant <= "01111110";
    type_cast_10310_wire_constant <= "01011101";
    type_cast_10312_wire_constant <= "01100100";
    type_cast_10320_wire_constant <= "01110011";
    type_cast_10322_wire_constant <= "00011001";
    type_cast_10330_wire_constant <= "10000001";
    type_cast_10332_wire_constant <= "01100000";
    type_cast_10340_wire_constant <= "11011100";
    type_cast_10342_wire_constant <= "01001111";
    type_cast_10350_wire_constant <= "00101010";
    type_cast_10352_wire_constant <= "00100010";
    type_cast_10360_wire_constant <= "10001000";
    type_cast_10362_wire_constant <= "10010000";
    type_cast_10370_wire_constant <= "11101110";
    type_cast_10372_wire_constant <= "01000110";
    type_cast_10380_wire_constant <= "00010100";
    type_cast_10382_wire_constant <= "10111000";
    type_cast_10390_wire_constant <= "01011110";
    type_cast_10392_wire_constant <= "11011110";
    type_cast_10400_wire_constant <= "11011011";
    type_cast_10402_wire_constant <= "00001011";
    type_cast_10410_wire_constant <= "00110010";
    type_cast_10412_wire_constant <= "11100000";
    type_cast_10420_wire_constant <= "00001010";
    type_cast_10422_wire_constant <= "00111010";
    type_cast_10430_wire_constant <= "00000110";
    type_cast_10432_wire_constant <= "01001001";
    type_cast_10440_wire_constant <= "01011100";
    type_cast_10442_wire_constant <= "00100100";
    type_cast_10450_wire_constant <= "11010011";
    type_cast_10452_wire_constant <= "11000010";
    type_cast_10460_wire_constant <= "01100010";
    type_cast_10462_wire_constant <= "10101100";
    type_cast_10470_wire_constant <= "10010101";
    type_cast_10472_wire_constant <= "10010001";
    type_cast_10480_wire_constant <= "01111001";
    type_cast_10482_wire_constant <= "11100100";
    type_cast_10490_wire_constant <= "11001000";
    type_cast_10492_wire_constant <= "11100111";
    type_cast_10500_wire_constant <= "01101101";
    type_cast_10502_wire_constant <= "00110111";
    type_cast_10510_wire_constant <= "11010101";
    type_cast_10512_wire_constant <= "10001101";
    type_cast_10520_wire_constant <= "10101001";
    type_cast_10522_wire_constant <= "01001110";
    type_cast_10530_wire_constant <= "01010110";
    type_cast_10532_wire_constant <= "01101100";
    type_cast_10540_wire_constant <= "11101010";
    type_cast_10542_wire_constant <= "11110100";
    type_cast_10550_wire_constant <= "01111010";
    type_cast_10552_wire_constant <= "01100101";
    type_cast_10560_wire_constant <= "00001000";
    type_cast_10562_wire_constant <= "10101110";
    type_cast_10570_wire_constant <= "01111000";
    type_cast_10572_wire_constant <= "10111010";
    type_cast_10580_wire_constant <= "00101110";
    type_cast_10582_wire_constant <= "00100101";
    type_cast_10590_wire_constant <= "10100110";
    type_cast_10592_wire_constant <= "00011100";
    type_cast_10600_wire_constant <= "11000110";
    type_cast_10602_wire_constant <= "10110100";
    type_cast_10610_wire_constant <= "11011101";
    type_cast_10612_wire_constant <= "11101000";
    type_cast_10620_wire_constant <= "00011111";
    type_cast_10622_wire_constant <= "01110100";
    type_cast_10630_wire_constant <= "10111101";
    type_cast_10632_wire_constant <= "01001011";
    type_cast_10640_wire_constant <= "10001010";
    type_cast_10642_wire_constant <= "10001011";
    type_cast_10650_wire_constant <= "00111110";
    type_cast_10652_wire_constant <= "01110000";
    type_cast_10660_wire_constant <= "01100110";
    type_cast_10662_wire_constant <= "10110101";
    type_cast_10670_wire_constant <= "00000011";
    type_cast_10672_wire_constant <= "01001000";
    type_cast_10680_wire_constant <= "00001110";
    type_cast_10682_wire_constant <= "11110110";
    type_cast_10690_wire_constant <= "00110101";
    type_cast_10692_wire_constant <= "01100001";
    type_cast_10700_wire_constant <= "10111001";
    type_cast_10702_wire_constant <= "01010111";
    type_cast_10710_wire_constant <= "11000001";
    type_cast_10712_wire_constant <= "10000110";
    type_cast_10720_wire_constant <= "10011110";
    type_cast_10722_wire_constant <= "00011101";
    type_cast_10730_wire_constant <= "11111000";
    type_cast_10732_wire_constant <= "11100001";
    type_cast_10740_wire_constant <= "00010001";
    type_cast_10742_wire_constant <= "10011000";
    type_cast_10750_wire_constant <= "11011001";
    type_cast_10752_wire_constant <= "01101001";
    type_cast_10760_wire_constant <= "10010100";
    type_cast_10762_wire_constant <= "10001110";
    type_cast_10770_wire_constant <= "00011110";
    type_cast_10772_wire_constant <= "10011011";
    type_cast_10780_wire_constant <= "11101001";
    type_cast_10782_wire_constant <= "10000111";
    type_cast_10790_wire_constant <= "01010101";
    type_cast_10792_wire_constant <= "11001110";
    type_cast_10800_wire_constant <= "11011111";
    type_cast_10802_wire_constant <= "00101000";
    type_cast_10810_wire_constant <= "10100001";
    type_cast_10812_wire_constant <= "10001100";
    type_cast_10820_wire_constant <= "00001101";
    type_cast_10822_wire_constant <= "10001001";
    type_cast_10830_wire_constant <= "11100110";
    type_cast_10832_wire_constant <= "10111111";
    type_cast_10840_wire_constant <= "01101000";
    type_cast_10842_wire_constant <= "01000010";
    type_cast_10850_wire_constant <= "10011001";
    type_cast_10852_wire_constant <= "01000001";
    type_cast_10860_wire_constant <= "00001111";
    type_cast_10862_wire_constant <= "00101101";
    type_cast_10870_wire_constant <= "01010100";
    type_cast_10872_wire_constant <= "10110000";
    type_cast_10880_wire_constant <= "00010110";
    type_cast_10882_wire_constant <= "10111011";
    type_cast_9610_wire_constant <= "01111100";
    type_cast_9612_wire_constant <= "01100011";
    type_cast_9620_wire_constant <= "01111011";
    type_cast_9622_wire_constant <= "01110111";
    type_cast_9630_wire_constant <= "01101011";
    type_cast_9632_wire_constant <= "11110010";
    type_cast_9640_wire_constant <= "11000101";
    type_cast_9642_wire_constant <= "01101111";
    type_cast_9650_wire_constant <= "00000001";
    type_cast_9652_wire_constant <= "00110000";
    type_cast_9660_wire_constant <= "00101011";
    type_cast_9662_wire_constant <= "01100111";
    type_cast_9670_wire_constant <= "11010111";
    type_cast_9672_wire_constant <= "11111110";
    type_cast_9680_wire_constant <= "01110110";
    type_cast_9682_wire_constant <= "10101011";
    type_cast_9690_wire_constant <= "10000010";
    type_cast_9692_wire_constant <= "11001010";
    type_cast_9700_wire_constant <= "01111101";
    type_cast_9702_wire_constant <= "11001001";
    type_cast_9710_wire_constant <= "01011001";
    type_cast_9712_wire_constant <= "11111010";
    type_cast_9720_wire_constant <= "11110000";
    type_cast_9722_wire_constant <= "01000111";
    type_cast_9730_wire_constant <= "11010100";
    type_cast_9732_wire_constant <= "10101101";
    type_cast_9740_wire_constant <= "10101111";
    type_cast_9742_wire_constant <= "10100010";
    type_cast_9750_wire_constant <= "10100100";
    type_cast_9752_wire_constant <= "10011100";
    type_cast_9760_wire_constant <= "11000000";
    type_cast_9762_wire_constant <= "01110010";
    type_cast_9770_wire_constant <= "11111101";
    type_cast_9772_wire_constant <= "10110111";
    type_cast_9780_wire_constant <= "00100110";
    type_cast_9782_wire_constant <= "10010011";
    type_cast_9790_wire_constant <= "00111111";
    type_cast_9792_wire_constant <= "00110110";
    type_cast_9800_wire_constant <= "11001100";
    type_cast_9802_wire_constant <= "11110111";
    type_cast_9810_wire_constant <= "10100101";
    type_cast_9812_wire_constant <= "00110100";
    type_cast_9820_wire_constant <= "11110001";
    type_cast_9822_wire_constant <= "11100101";
    type_cast_9830_wire_constant <= "11011000";
    type_cast_9832_wire_constant <= "01110001";
    type_cast_9840_wire_constant <= "00010101";
    type_cast_9842_wire_constant <= "00110001";
    type_cast_9850_wire_constant <= "11000111";
    type_cast_9852_wire_constant <= "00000100";
    type_cast_9860_wire_constant <= "11000011";
    type_cast_9862_wire_constant <= "00100011";
    type_cast_9870_wire_constant <= "10010110";
    type_cast_9872_wire_constant <= "00011000";
    type_cast_9880_wire_constant <= "10011010";
    type_cast_9882_wire_constant <= "00000101";
    type_cast_9890_wire_constant <= "00010010";
    type_cast_9892_wire_constant <= "00000111";
    type_cast_9900_wire_constant <= "11100010";
    type_cast_9902_wire_constant <= "10000000";
    type_cast_9910_wire_constant <= "00100111";
    type_cast_9912_wire_constant <= "11101011";
    type_cast_9920_wire_constant <= "01110101";
    type_cast_9922_wire_constant <= "10110010";
    type_cast_9930_wire_constant <= "10000011";
    type_cast_9932_wire_constant <= "00001001";
    type_cast_9940_wire_constant <= "00011010";
    type_cast_9942_wire_constant <= "00101100";
    type_cast_9950_wire_constant <= "01101110";
    type_cast_9952_wire_constant <= "00011011";
    type_cast_9960_wire_constant <= "10100000";
    type_cast_9962_wire_constant <= "01011010";
    type_cast_9970_wire_constant <= "00111011";
    type_cast_9972_wire_constant <= "01010010";
    type_cast_9980_wire_constant <= "10110011";
    type_cast_9982_wire_constant <= "11010110";
    type_cast_9990_wire_constant <= "11100011";
    type_cast_9992_wire_constant <= "00101001";
    -- flow-through select operator MUX_10003_inst
    MA39_10004 <= type_cast_10000_wire_constant when (BITSEL_u8_u1_9998_wire(0) /=  '0') else type_cast_10002_wire_constant;
    -- flow-through select operator MUX_10013_inst
    MA40_10014 <= type_cast_10010_wire_constant when (BITSEL_u8_u1_10008_wire(0) /=  '0') else type_cast_10012_wire_constant;
    -- flow-through select operator MUX_10023_inst
    MA41_10024 <= type_cast_10020_wire_constant when (BITSEL_u8_u1_10018_wire(0) /=  '0') else type_cast_10022_wire_constant;
    -- flow-through select operator MUX_10033_inst
    MA42_10034 <= type_cast_10030_wire_constant when (BITSEL_u8_u1_10028_wire(0) /=  '0') else type_cast_10032_wire_constant;
    -- flow-through select operator MUX_10043_inst
    MA43_10044 <= type_cast_10040_wire_constant when (BITSEL_u8_u1_10038_wire(0) /=  '0') else type_cast_10042_wire_constant;
    -- flow-through select operator MUX_10053_inst
    MA44_10054 <= type_cast_10050_wire_constant when (BITSEL_u8_u1_10048_wire(0) /=  '0') else type_cast_10052_wire_constant;
    -- flow-through select operator MUX_10063_inst
    MA45_10064 <= type_cast_10060_wire_constant when (BITSEL_u8_u1_10058_wire(0) /=  '0') else type_cast_10062_wire_constant;
    -- flow-through select operator MUX_10073_inst
    MA46_10074 <= type_cast_10070_wire_constant when (BITSEL_u8_u1_10068_wire(0) /=  '0') else type_cast_10072_wire_constant;
    -- flow-through select operator MUX_10083_inst
    MA47_10084 <= type_cast_10080_wire_constant when (BITSEL_u8_u1_10078_wire(0) /=  '0') else type_cast_10082_wire_constant;
    -- flow-through select operator MUX_10093_inst
    MA48_10094 <= type_cast_10090_wire_constant when (BITSEL_u8_u1_10088_wire(0) /=  '0') else type_cast_10092_wire_constant;
    -- flow-through select operator MUX_10103_inst
    MA49_10104 <= type_cast_10100_wire_constant when (BITSEL_u8_u1_10098_wire(0) /=  '0') else type_cast_10102_wire_constant;
    -- flow-through select operator MUX_10113_inst
    MA50_10114 <= type_cast_10110_wire_constant when (BITSEL_u8_u1_10108_wire(0) /=  '0') else type_cast_10112_wire_constant;
    -- flow-through select operator MUX_10123_inst
    MA51_10124 <= type_cast_10120_wire_constant when (BITSEL_u8_u1_10118_wire(0) /=  '0') else type_cast_10122_wire_constant;
    -- flow-through select operator MUX_10133_inst
    MA52_10134 <= type_cast_10130_wire_constant when (BITSEL_u8_u1_10128_wire(0) /=  '0') else type_cast_10132_wire_constant;
    -- flow-through select operator MUX_10143_inst
    MA53_10144 <= type_cast_10140_wire_constant when (BITSEL_u8_u1_10138_wire(0) /=  '0') else type_cast_10142_wire_constant;
    -- flow-through select operator MUX_10153_inst
    MA54_10154 <= type_cast_10150_wire_constant when (BITSEL_u8_u1_10148_wire(0) /=  '0') else type_cast_10152_wire_constant;
    -- flow-through select operator MUX_10163_inst
    MA55_10164 <= type_cast_10160_wire_constant when (BITSEL_u8_u1_10158_wire(0) /=  '0') else type_cast_10162_wire_constant;
    -- flow-through select operator MUX_10173_inst
    MA56_10174 <= type_cast_10170_wire_constant when (BITSEL_u8_u1_10168_wire(0) /=  '0') else type_cast_10172_wire_constant;
    -- flow-through select operator MUX_10183_inst
    MA57_10184 <= type_cast_10180_wire_constant when (BITSEL_u8_u1_10178_wire(0) /=  '0') else type_cast_10182_wire_constant;
    -- flow-through select operator MUX_10193_inst
    MA58_10194 <= type_cast_10190_wire_constant when (BITSEL_u8_u1_10188_wire(0) /=  '0') else type_cast_10192_wire_constant;
    -- flow-through select operator MUX_10203_inst
    MA59_10204 <= type_cast_10200_wire_constant when (BITSEL_u8_u1_10198_wire(0) /=  '0') else type_cast_10202_wire_constant;
    -- flow-through select operator MUX_10213_inst
    MA60_10214 <= type_cast_10210_wire_constant when (BITSEL_u8_u1_10208_wire(0) /=  '0') else type_cast_10212_wire_constant;
    -- flow-through select operator MUX_10223_inst
    MA61_10224 <= type_cast_10220_wire_constant when (BITSEL_u8_u1_10218_wire(0) /=  '0') else type_cast_10222_wire_constant;
    -- flow-through select operator MUX_10233_inst
    MA62_10234 <= type_cast_10230_wire_constant when (BITSEL_u8_u1_10228_wire(0) /=  '0') else type_cast_10232_wire_constant;
    -- flow-through select operator MUX_10243_inst
    MA63_10244 <= type_cast_10240_wire_constant when (BITSEL_u8_u1_10238_wire(0) /=  '0') else type_cast_10242_wire_constant;
    -- flow-through select operator MUX_10253_inst
    MA64_10254 <= type_cast_10250_wire_constant when (BITSEL_u8_u1_10248_wire(0) /=  '0') else type_cast_10252_wire_constant;
    -- flow-through select operator MUX_10263_inst
    MA65_10264 <= type_cast_10260_wire_constant when (BITSEL_u8_u1_10258_wire(0) /=  '0') else type_cast_10262_wire_constant;
    -- flow-through select operator MUX_10273_inst
    MA66_10274 <= type_cast_10270_wire_constant when (BITSEL_u8_u1_10268_wire(0) /=  '0') else type_cast_10272_wire_constant;
    -- flow-through select operator MUX_10283_inst
    MA67_10284 <= type_cast_10280_wire_constant when (BITSEL_u8_u1_10278_wire(0) /=  '0') else type_cast_10282_wire_constant;
    -- flow-through select operator MUX_10293_inst
    MA68_10294 <= type_cast_10290_wire_constant when (BITSEL_u8_u1_10288_wire(0) /=  '0') else type_cast_10292_wire_constant;
    -- flow-through select operator MUX_10303_inst
    MA69_10304 <= type_cast_10300_wire_constant when (BITSEL_u8_u1_10298_wire(0) /=  '0') else type_cast_10302_wire_constant;
    -- flow-through select operator MUX_10313_inst
    MA70_10314 <= type_cast_10310_wire_constant when (BITSEL_u8_u1_10308_wire(0) /=  '0') else type_cast_10312_wire_constant;
    -- flow-through select operator MUX_10323_inst
    MA71_10324 <= type_cast_10320_wire_constant when (BITSEL_u8_u1_10318_wire(0) /=  '0') else type_cast_10322_wire_constant;
    -- flow-through select operator MUX_10333_inst
    MA72_10334 <= type_cast_10330_wire_constant when (BITSEL_u8_u1_10328_wire(0) /=  '0') else type_cast_10332_wire_constant;
    -- flow-through select operator MUX_10343_inst
    MA73_10344 <= type_cast_10340_wire_constant when (BITSEL_u8_u1_10338_wire(0) /=  '0') else type_cast_10342_wire_constant;
    -- flow-through select operator MUX_10353_inst
    MA74_10354 <= type_cast_10350_wire_constant when (BITSEL_u8_u1_10348_wire(0) /=  '0') else type_cast_10352_wire_constant;
    -- flow-through select operator MUX_10363_inst
    MA75_10364 <= type_cast_10360_wire_constant when (BITSEL_u8_u1_10358_wire(0) /=  '0') else type_cast_10362_wire_constant;
    -- flow-through select operator MUX_10373_inst
    MA76_10374 <= type_cast_10370_wire_constant when (BITSEL_u8_u1_10368_wire(0) /=  '0') else type_cast_10372_wire_constant;
    -- flow-through select operator MUX_10383_inst
    MA77_10384 <= type_cast_10380_wire_constant when (BITSEL_u8_u1_10378_wire(0) /=  '0') else type_cast_10382_wire_constant;
    -- flow-through select operator MUX_10393_inst
    MA78_10394 <= type_cast_10390_wire_constant when (BITSEL_u8_u1_10388_wire(0) /=  '0') else type_cast_10392_wire_constant;
    -- flow-through select operator MUX_10403_inst
    MA79_10404 <= type_cast_10400_wire_constant when (BITSEL_u8_u1_10398_wire(0) /=  '0') else type_cast_10402_wire_constant;
    -- flow-through select operator MUX_10413_inst
    MA80_10414 <= type_cast_10410_wire_constant when (BITSEL_u8_u1_10408_wire(0) /=  '0') else type_cast_10412_wire_constant;
    -- flow-through select operator MUX_10423_inst
    MA81_10424 <= type_cast_10420_wire_constant when (BITSEL_u8_u1_10418_wire(0) /=  '0') else type_cast_10422_wire_constant;
    -- flow-through select operator MUX_10433_inst
    MA82_10434 <= type_cast_10430_wire_constant when (BITSEL_u8_u1_10428_wire(0) /=  '0') else type_cast_10432_wire_constant;
    -- flow-through select operator MUX_10443_inst
    MA83_10444 <= type_cast_10440_wire_constant when (BITSEL_u8_u1_10438_wire(0) /=  '0') else type_cast_10442_wire_constant;
    -- flow-through select operator MUX_10453_inst
    MA84_10454 <= type_cast_10450_wire_constant when (BITSEL_u8_u1_10448_wire(0) /=  '0') else type_cast_10452_wire_constant;
    -- flow-through select operator MUX_10463_inst
    MA85_10464 <= type_cast_10460_wire_constant when (BITSEL_u8_u1_10458_wire(0) /=  '0') else type_cast_10462_wire_constant;
    -- flow-through select operator MUX_10473_inst
    MA86_10474 <= type_cast_10470_wire_constant when (BITSEL_u8_u1_10468_wire(0) /=  '0') else type_cast_10472_wire_constant;
    -- flow-through select operator MUX_10483_inst
    MA87_10484 <= type_cast_10480_wire_constant when (BITSEL_u8_u1_10478_wire(0) /=  '0') else type_cast_10482_wire_constant;
    -- flow-through select operator MUX_10493_inst
    MA88_10494 <= type_cast_10490_wire_constant when (BITSEL_u8_u1_10488_wire(0) /=  '0') else type_cast_10492_wire_constant;
    -- flow-through select operator MUX_10503_inst
    MA89_10504 <= type_cast_10500_wire_constant when (BITSEL_u8_u1_10498_wire(0) /=  '0') else type_cast_10502_wire_constant;
    -- flow-through select operator MUX_10513_inst
    MA90_10514 <= type_cast_10510_wire_constant when (BITSEL_u8_u1_10508_wire(0) /=  '0') else type_cast_10512_wire_constant;
    -- flow-through select operator MUX_10523_inst
    MA91_10524 <= type_cast_10520_wire_constant when (BITSEL_u8_u1_10518_wire(0) /=  '0') else type_cast_10522_wire_constant;
    -- flow-through select operator MUX_10533_inst
    MA92_10534 <= type_cast_10530_wire_constant when (BITSEL_u8_u1_10528_wire(0) /=  '0') else type_cast_10532_wire_constant;
    -- flow-through select operator MUX_10543_inst
    MA93_10544 <= type_cast_10540_wire_constant when (BITSEL_u8_u1_10538_wire(0) /=  '0') else type_cast_10542_wire_constant;
    -- flow-through select operator MUX_10553_inst
    MA94_10554 <= type_cast_10550_wire_constant when (BITSEL_u8_u1_10548_wire(0) /=  '0') else type_cast_10552_wire_constant;
    -- flow-through select operator MUX_10563_inst
    MA95_10564 <= type_cast_10560_wire_constant when (BITSEL_u8_u1_10558_wire(0) /=  '0') else type_cast_10562_wire_constant;
    -- flow-through select operator MUX_10573_inst
    MA96_10574 <= type_cast_10570_wire_constant when (BITSEL_u8_u1_10568_wire(0) /=  '0') else type_cast_10572_wire_constant;
    -- flow-through select operator MUX_10583_inst
    MA97_10584 <= type_cast_10580_wire_constant when (BITSEL_u8_u1_10578_wire(0) /=  '0') else type_cast_10582_wire_constant;
    -- flow-through select operator MUX_10593_inst
    MA98_10594 <= type_cast_10590_wire_constant when (BITSEL_u8_u1_10588_wire(0) /=  '0') else type_cast_10592_wire_constant;
    -- flow-through select operator MUX_10603_inst
    MA99_10604 <= type_cast_10600_wire_constant when (BITSEL_u8_u1_10598_wire(0) /=  '0') else type_cast_10602_wire_constant;
    -- flow-through select operator MUX_10613_inst
    MA100_10614 <= type_cast_10610_wire_constant when (BITSEL_u8_u1_10608_wire(0) /=  '0') else type_cast_10612_wire_constant;
    -- flow-through select operator MUX_10623_inst
    MA101_10624 <= type_cast_10620_wire_constant when (BITSEL_u8_u1_10618_wire(0) /=  '0') else type_cast_10622_wire_constant;
    -- flow-through select operator MUX_10633_inst
    MA102_10634 <= type_cast_10630_wire_constant when (BITSEL_u8_u1_10628_wire(0) /=  '0') else type_cast_10632_wire_constant;
    -- flow-through select operator MUX_10643_inst
    MA103_10644 <= type_cast_10640_wire_constant when (BITSEL_u8_u1_10638_wire(0) /=  '0') else type_cast_10642_wire_constant;
    -- flow-through select operator MUX_10653_inst
    MA104_10654 <= type_cast_10650_wire_constant when (BITSEL_u8_u1_10648_wire(0) /=  '0') else type_cast_10652_wire_constant;
    -- flow-through select operator MUX_10663_inst
    MA105_10664 <= type_cast_10660_wire_constant when (BITSEL_u8_u1_10658_wire(0) /=  '0') else type_cast_10662_wire_constant;
    -- flow-through select operator MUX_10673_inst
    MA106_10674 <= type_cast_10670_wire_constant when (BITSEL_u8_u1_10668_wire(0) /=  '0') else type_cast_10672_wire_constant;
    -- flow-through select operator MUX_10683_inst
    MA107_10684 <= type_cast_10680_wire_constant when (BITSEL_u8_u1_10678_wire(0) /=  '0') else type_cast_10682_wire_constant;
    -- flow-through select operator MUX_10693_inst
    MA108_10694 <= type_cast_10690_wire_constant when (BITSEL_u8_u1_10688_wire(0) /=  '0') else type_cast_10692_wire_constant;
    -- flow-through select operator MUX_10703_inst
    MA109_10704 <= type_cast_10700_wire_constant when (BITSEL_u8_u1_10698_wire(0) /=  '0') else type_cast_10702_wire_constant;
    -- flow-through select operator MUX_10713_inst
    MA110_10714 <= type_cast_10710_wire_constant when (BITSEL_u8_u1_10708_wire(0) /=  '0') else type_cast_10712_wire_constant;
    -- flow-through select operator MUX_10723_inst
    MA111_10724 <= type_cast_10720_wire_constant when (BITSEL_u8_u1_10718_wire(0) /=  '0') else type_cast_10722_wire_constant;
    -- flow-through select operator MUX_10733_inst
    MA112_10734 <= type_cast_10730_wire_constant when (BITSEL_u8_u1_10728_wire(0) /=  '0') else type_cast_10732_wire_constant;
    -- flow-through select operator MUX_10743_inst
    MA113_10744 <= type_cast_10740_wire_constant when (BITSEL_u8_u1_10738_wire(0) /=  '0') else type_cast_10742_wire_constant;
    -- flow-through select operator MUX_10753_inst
    MA114_10754 <= type_cast_10750_wire_constant when (BITSEL_u8_u1_10748_wire(0) /=  '0') else type_cast_10752_wire_constant;
    -- flow-through select operator MUX_10763_inst
    MA115_10764 <= type_cast_10760_wire_constant when (BITSEL_u8_u1_10758_wire(0) /=  '0') else type_cast_10762_wire_constant;
    -- flow-through select operator MUX_10773_inst
    MA116_10774 <= type_cast_10770_wire_constant when (BITSEL_u8_u1_10768_wire(0) /=  '0') else type_cast_10772_wire_constant;
    -- flow-through select operator MUX_10783_inst
    MA117_10784 <= type_cast_10780_wire_constant when (BITSEL_u8_u1_10778_wire(0) /=  '0') else type_cast_10782_wire_constant;
    -- flow-through select operator MUX_10793_inst
    MA118_10794 <= type_cast_10790_wire_constant when (BITSEL_u8_u1_10788_wire(0) /=  '0') else type_cast_10792_wire_constant;
    -- flow-through select operator MUX_10803_inst
    MA119_10804 <= type_cast_10800_wire_constant when (BITSEL_u8_u1_10798_wire(0) /=  '0') else type_cast_10802_wire_constant;
    -- flow-through select operator MUX_10813_inst
    MA120_10814 <= type_cast_10810_wire_constant when (BITSEL_u8_u1_10808_wire(0) /=  '0') else type_cast_10812_wire_constant;
    -- flow-through select operator MUX_10823_inst
    MA121_10824 <= type_cast_10820_wire_constant when (BITSEL_u8_u1_10818_wire(0) /=  '0') else type_cast_10822_wire_constant;
    -- flow-through select operator MUX_10833_inst
    MA122_10834 <= type_cast_10830_wire_constant when (BITSEL_u8_u1_10828_wire(0) /=  '0') else type_cast_10832_wire_constant;
    -- flow-through select operator MUX_10843_inst
    MA123_10844 <= type_cast_10840_wire_constant when (BITSEL_u8_u1_10838_wire(0) /=  '0') else type_cast_10842_wire_constant;
    -- flow-through select operator MUX_10853_inst
    MA124_10854 <= type_cast_10850_wire_constant when (BITSEL_u8_u1_10848_wire(0) /=  '0') else type_cast_10852_wire_constant;
    -- flow-through select operator MUX_10863_inst
    MA125_10864 <= type_cast_10860_wire_constant when (BITSEL_u8_u1_10858_wire(0) /=  '0') else type_cast_10862_wire_constant;
    -- flow-through select operator MUX_10873_inst
    MA126_10874 <= type_cast_10870_wire_constant when (BITSEL_u8_u1_10868_wire(0) /=  '0') else type_cast_10872_wire_constant;
    -- flow-through select operator MUX_10883_inst
    MA127_10884 <= type_cast_10880_wire_constant when (BITSEL_u8_u1_10878_wire(0) /=  '0') else type_cast_10882_wire_constant;
    -- flow-through select operator MUX_10891_inst
    MB0_10892 <= MA1_9624 when (BITSEL_u8_u1_10888_wire(0) /=  '0') else MA0_9614;
    -- flow-through select operator MUX_10899_inst
    MB1_10900 <= MA3_9644 when (BITSEL_u8_u1_10896_wire(0) /=  '0') else MA2_9634;
    -- flow-through select operator MUX_10907_inst
    MB2_10908 <= MA5_9664 when (BITSEL_u8_u1_10904_wire(0) /=  '0') else MA4_9654;
    -- flow-through select operator MUX_10915_inst
    MB3_10916 <= MA7_9684 when (BITSEL_u8_u1_10912_wire(0) /=  '0') else MA6_9674;
    -- flow-through select operator MUX_10923_inst
    MB4_10924 <= MA9_9704 when (BITSEL_u8_u1_10920_wire(0) /=  '0') else MA8_9694;
    -- flow-through select operator MUX_10931_inst
    MB5_10932 <= MA11_9724 when (BITSEL_u8_u1_10928_wire(0) /=  '0') else MA10_9714;
    -- flow-through select operator MUX_10939_inst
    MB6_10940 <= MA13_9744 when (BITSEL_u8_u1_10936_wire(0) /=  '0') else MA12_9734;
    -- flow-through select operator MUX_10947_inst
    MB7_10948 <= MA15_9764 when (BITSEL_u8_u1_10944_wire(0) /=  '0') else MA14_9754;
    -- flow-through select operator MUX_10955_inst
    MB8_10956 <= MA17_9784 when (BITSEL_u8_u1_10952_wire(0) /=  '0') else MA16_9774;
    -- flow-through select operator MUX_10963_inst
    MB9_10964 <= MA19_9804 when (BITSEL_u8_u1_10960_wire(0) /=  '0') else MA18_9794;
    -- flow-through select operator MUX_10971_inst
    MB10_10972 <= MA21_9824 when (BITSEL_u8_u1_10968_wire(0) /=  '0') else MA20_9814;
    -- flow-through select operator MUX_10979_inst
    MB11_10980 <= MA23_9844 when (BITSEL_u8_u1_10976_wire(0) /=  '0') else MA22_9834;
    -- flow-through select operator MUX_10987_inst
    MB12_10988 <= MA25_9864 when (BITSEL_u8_u1_10984_wire(0) /=  '0') else MA24_9854;
    -- flow-through select operator MUX_10995_inst
    MB13_10996 <= MA27_9884 when (BITSEL_u8_u1_10992_wire(0) /=  '0') else MA26_9874;
    -- flow-through select operator MUX_11003_inst
    MB14_11004 <= MA29_9904 when (BITSEL_u8_u1_11000_wire(0) /=  '0') else MA28_9894;
    -- flow-through select operator MUX_11011_inst
    MB15_11012 <= MA31_9924 when (BITSEL_u8_u1_11008_wire(0) /=  '0') else MA30_9914;
    -- flow-through select operator MUX_11019_inst
    MB16_11020 <= MA33_9944 when (BITSEL_u8_u1_11016_wire(0) /=  '0') else MA32_9934;
    -- flow-through select operator MUX_11027_inst
    MB17_11028 <= MA35_9964 when (BITSEL_u8_u1_11024_wire(0) /=  '0') else MA34_9954;
    -- flow-through select operator MUX_11035_inst
    MB18_11036 <= MA37_9984 when (BITSEL_u8_u1_11032_wire(0) /=  '0') else MA36_9974;
    -- flow-through select operator MUX_11043_inst
    MB19_11044 <= MA39_10004 when (BITSEL_u8_u1_11040_wire(0) /=  '0') else MA38_9994;
    -- flow-through select operator MUX_11051_inst
    MB20_11052 <= MA41_10024 when (BITSEL_u8_u1_11048_wire(0) /=  '0') else MA40_10014;
    -- flow-through select operator MUX_11059_inst
    MB21_11060 <= MA43_10044 when (BITSEL_u8_u1_11056_wire(0) /=  '0') else MA42_10034;
    -- flow-through select operator MUX_11067_inst
    MB22_11068 <= MA45_10064 when (BITSEL_u8_u1_11064_wire(0) /=  '0') else MA44_10054;
    -- flow-through select operator MUX_11075_inst
    MB23_11076 <= MA47_10084 when (BITSEL_u8_u1_11072_wire(0) /=  '0') else MA46_10074;
    -- flow-through select operator MUX_11083_inst
    MB24_11084 <= MA49_10104 when (BITSEL_u8_u1_11080_wire(0) /=  '0') else MA48_10094;
    -- flow-through select operator MUX_11091_inst
    MB25_11092 <= MA51_10124 when (BITSEL_u8_u1_11088_wire(0) /=  '0') else MA50_10114;
    -- flow-through select operator MUX_11099_inst
    MB26_11100 <= MA53_10144 when (BITSEL_u8_u1_11096_wire(0) /=  '0') else MA52_10134;
    -- flow-through select operator MUX_11107_inst
    MB27_11108 <= MA55_10164 when (BITSEL_u8_u1_11104_wire(0) /=  '0') else MA54_10154;
    -- flow-through select operator MUX_11115_inst
    MB28_11116 <= MA57_10184 when (BITSEL_u8_u1_11112_wire(0) /=  '0') else MA56_10174;
    -- flow-through select operator MUX_11123_inst
    MB29_11124 <= MA59_10204 when (BITSEL_u8_u1_11120_wire(0) /=  '0') else MA58_10194;
    -- flow-through select operator MUX_11131_inst
    MB30_11132 <= MA61_10224 when (BITSEL_u8_u1_11128_wire(0) /=  '0') else MA60_10214;
    -- flow-through select operator MUX_11139_inst
    MB31_11140 <= MA63_10244 when (BITSEL_u8_u1_11136_wire(0) /=  '0') else MA62_10234;
    -- flow-through select operator MUX_11147_inst
    MB32_11148 <= MA65_10264 when (BITSEL_u8_u1_11144_wire(0) /=  '0') else MA64_10254;
    -- flow-through select operator MUX_11155_inst
    MB33_11156 <= MA67_10284 when (BITSEL_u8_u1_11152_wire(0) /=  '0') else MA66_10274;
    -- flow-through select operator MUX_11163_inst
    MB34_11164 <= MA69_10304 when (BITSEL_u8_u1_11160_wire(0) /=  '0') else MA68_10294;
    -- flow-through select operator MUX_11171_inst
    MB35_11172 <= MA71_10324 when (BITSEL_u8_u1_11168_wire(0) /=  '0') else MA70_10314;
    -- flow-through select operator MUX_11179_inst
    MB36_11180 <= MA73_10344 when (BITSEL_u8_u1_11176_wire(0) /=  '0') else MA72_10334;
    -- flow-through select operator MUX_11187_inst
    MB37_11188 <= MA75_10364 when (BITSEL_u8_u1_11184_wire(0) /=  '0') else MA74_10354;
    -- flow-through select operator MUX_11195_inst
    MB38_11196 <= MA77_10384 when (BITSEL_u8_u1_11192_wire(0) /=  '0') else MA76_10374;
    -- flow-through select operator MUX_11203_inst
    MB39_11204 <= MA79_10404 when (BITSEL_u8_u1_11200_wire(0) /=  '0') else MA78_10394;
    -- flow-through select operator MUX_11211_inst
    MB40_11212 <= MA81_10424 when (BITSEL_u8_u1_11208_wire(0) /=  '0') else MA80_10414;
    -- flow-through select operator MUX_11219_inst
    MB41_11220 <= MA83_10444 when (BITSEL_u8_u1_11216_wire(0) /=  '0') else MA82_10434;
    -- flow-through select operator MUX_11227_inst
    MB42_11228 <= MA85_10464 when (BITSEL_u8_u1_11224_wire(0) /=  '0') else MA84_10454;
    -- flow-through select operator MUX_11235_inst
    MB43_11236 <= MA87_10484 when (BITSEL_u8_u1_11232_wire(0) /=  '0') else MA86_10474;
    -- flow-through select operator MUX_11243_inst
    MB44_11244 <= MA89_10504 when (BITSEL_u8_u1_11240_wire(0) /=  '0') else MA88_10494;
    -- flow-through select operator MUX_11251_inst
    MB45_11252 <= MA91_10524 when (BITSEL_u8_u1_11248_wire(0) /=  '0') else MA90_10514;
    -- flow-through select operator MUX_11259_inst
    MB46_11260 <= MA93_10544 when (BITSEL_u8_u1_11256_wire(0) /=  '0') else MA92_10534;
    -- flow-through select operator MUX_11267_inst
    MB47_11268 <= MA95_10564 when (BITSEL_u8_u1_11264_wire(0) /=  '0') else MA94_10554;
    -- flow-through select operator MUX_11275_inst
    MB48_11276 <= MA97_10584 when (BITSEL_u8_u1_11272_wire(0) /=  '0') else MA96_10574;
    -- flow-through select operator MUX_11283_inst
    MB49_11284 <= MA99_10604 when (BITSEL_u8_u1_11280_wire(0) /=  '0') else MA98_10594;
    -- flow-through select operator MUX_11291_inst
    MB50_11292 <= MA101_10624 when (BITSEL_u8_u1_11288_wire(0) /=  '0') else MA100_10614;
    -- flow-through select operator MUX_11299_inst
    MB51_11300 <= MA103_10644 when (BITSEL_u8_u1_11296_wire(0) /=  '0') else MA102_10634;
    -- flow-through select operator MUX_11307_inst
    MB52_11308 <= MA105_10664 when (BITSEL_u8_u1_11304_wire(0) /=  '0') else MA104_10654;
    -- flow-through select operator MUX_11315_inst
    MB53_11316 <= MA107_10684 when (BITSEL_u8_u1_11312_wire(0) /=  '0') else MA106_10674;
    -- flow-through select operator MUX_11323_inst
    MB54_11324 <= MA109_10704 when (BITSEL_u8_u1_11320_wire(0) /=  '0') else MA108_10694;
    -- flow-through select operator MUX_11331_inst
    MB55_11332 <= MA111_10724 when (BITSEL_u8_u1_11328_wire(0) /=  '0') else MA110_10714;
    -- flow-through select operator MUX_11339_inst
    MB56_11340 <= MA113_10744 when (BITSEL_u8_u1_11336_wire(0) /=  '0') else MA112_10734;
    -- flow-through select operator MUX_11347_inst
    MB57_11348 <= MA115_10764 when (BITSEL_u8_u1_11344_wire(0) /=  '0') else MA114_10754;
    -- flow-through select operator MUX_11355_inst
    MB58_11356 <= MA117_10784 when (BITSEL_u8_u1_11352_wire(0) /=  '0') else MA116_10774;
    -- flow-through select operator MUX_11363_inst
    MB59_11364 <= MA119_10804 when (BITSEL_u8_u1_11360_wire(0) /=  '0') else MA118_10794;
    -- flow-through select operator MUX_11371_inst
    MB60_11372 <= MA121_10824 when (BITSEL_u8_u1_11368_wire(0) /=  '0') else MA120_10814;
    -- flow-through select operator MUX_11379_inst
    MB61_11380 <= MA123_10844 when (BITSEL_u8_u1_11376_wire(0) /=  '0') else MA122_10834;
    -- flow-through select operator MUX_11387_inst
    MB62_11388 <= MA125_10864 when (BITSEL_u8_u1_11384_wire(0) /=  '0') else MA124_10854;
    -- flow-through select operator MUX_11395_inst
    MB63_11396 <= MA127_10884 when (BITSEL_u8_u1_11392_wire(0) /=  '0') else MA126_10874;
    -- flow-through select operator MUX_11403_inst
    MC0_11404 <= MB1_10900 when (BITSEL_u8_u1_11400_wire(0) /=  '0') else MB0_10892;
    -- flow-through select operator MUX_11411_inst
    MC1_11412 <= MB3_10916 when (BITSEL_u8_u1_11408_wire(0) /=  '0') else MB2_10908;
    -- flow-through select operator MUX_11419_inst
    MC2_11420 <= MB5_10932 when (BITSEL_u8_u1_11416_wire(0) /=  '0') else MB4_10924;
    -- flow-through select operator MUX_11427_inst
    MC3_11428 <= MB7_10948 when (BITSEL_u8_u1_11424_wire(0) /=  '0') else MB6_10940;
    -- flow-through select operator MUX_11435_inst
    MC4_11436 <= MB9_10964 when (BITSEL_u8_u1_11432_wire(0) /=  '0') else MB8_10956;
    -- flow-through select operator MUX_11443_inst
    MC5_11444 <= MB11_10980 when (BITSEL_u8_u1_11440_wire(0) /=  '0') else MB10_10972;
    -- flow-through select operator MUX_11451_inst
    MC6_11452 <= MB13_10996 when (BITSEL_u8_u1_11448_wire(0) /=  '0') else MB12_10988;
    -- flow-through select operator MUX_11459_inst
    MC7_11460 <= MB15_11012 when (BITSEL_u8_u1_11456_wire(0) /=  '0') else MB14_11004;
    -- flow-through select operator MUX_11467_inst
    MC8_11468 <= MB17_11028 when (BITSEL_u8_u1_11464_wire(0) /=  '0') else MB16_11020;
    -- flow-through select operator MUX_11475_inst
    MC9_11476 <= MB19_11044 when (BITSEL_u8_u1_11472_wire(0) /=  '0') else MB18_11036;
    -- flow-through select operator MUX_11483_inst
    MC10_11484 <= MB21_11060 when (BITSEL_u8_u1_11480_wire(0) /=  '0') else MB20_11052;
    -- flow-through select operator MUX_11491_inst
    MC11_11492 <= MB23_11076 when (BITSEL_u8_u1_11488_wire(0) /=  '0') else MB22_11068;
    -- flow-through select operator MUX_11499_inst
    MC12_11500 <= MB25_11092 when (BITSEL_u8_u1_11496_wire(0) /=  '0') else MB24_11084;
    -- flow-through select operator MUX_11507_inst
    MC13_11508 <= MB27_11108 when (BITSEL_u8_u1_11504_wire(0) /=  '0') else MB26_11100;
    -- flow-through select operator MUX_11515_inst
    MC14_11516 <= MB29_11124 when (BITSEL_u8_u1_11512_wire(0) /=  '0') else MB28_11116;
    -- flow-through select operator MUX_11523_inst
    MC15_11524 <= MB31_11140 when (BITSEL_u8_u1_11520_wire(0) /=  '0') else MB30_11132;
    -- flow-through select operator MUX_11531_inst
    MC16_11532 <= MB33_11156 when (BITSEL_u8_u1_11528_wire(0) /=  '0') else MB32_11148;
    -- flow-through select operator MUX_11539_inst
    MC17_11540 <= MB35_11172 when (BITSEL_u8_u1_11536_wire(0) /=  '0') else MB34_11164;
    -- flow-through select operator MUX_11547_inst
    MC18_11548 <= MB37_11188 when (BITSEL_u8_u1_11544_wire(0) /=  '0') else MB36_11180;
    -- flow-through select operator MUX_11555_inst
    MC19_11556 <= MB39_11204 when (BITSEL_u8_u1_11552_wire(0) /=  '0') else MB38_11196;
    -- flow-through select operator MUX_11563_inst
    MC20_11564 <= MB41_11220 when (BITSEL_u8_u1_11560_wire(0) /=  '0') else MB40_11212;
    -- flow-through select operator MUX_11571_inst
    MC21_11572 <= MB43_11236 when (BITSEL_u8_u1_11568_wire(0) /=  '0') else MB42_11228;
    -- flow-through select operator MUX_11579_inst
    MC22_11580 <= MB45_11252 when (BITSEL_u8_u1_11576_wire(0) /=  '0') else MB44_11244;
    -- flow-through select operator MUX_11587_inst
    MC23_11588 <= MB47_11268 when (BITSEL_u8_u1_11584_wire(0) /=  '0') else MB46_11260;
    -- flow-through select operator MUX_11595_inst
    MC24_11596 <= MB49_11284 when (BITSEL_u8_u1_11592_wire(0) /=  '0') else MB48_11276;
    -- flow-through select operator MUX_11603_inst
    MC25_11604 <= MB51_11300 when (BITSEL_u8_u1_11600_wire(0) /=  '0') else MB50_11292;
    -- flow-through select operator MUX_11611_inst
    MC26_11612 <= MB53_11316 when (BITSEL_u8_u1_11608_wire(0) /=  '0') else MB52_11308;
    -- flow-through select operator MUX_11619_inst
    MC27_11620 <= MB55_11332 when (BITSEL_u8_u1_11616_wire(0) /=  '0') else MB54_11324;
    -- flow-through select operator MUX_11627_inst
    MC28_11628 <= MB57_11348 when (BITSEL_u8_u1_11624_wire(0) /=  '0') else MB56_11340;
    -- flow-through select operator MUX_11635_inst
    MC29_11636 <= MB59_11364 when (BITSEL_u8_u1_11632_wire(0) /=  '0') else MB58_11356;
    -- flow-through select operator MUX_11643_inst
    MC30_11644 <= MB61_11380 when (BITSEL_u8_u1_11640_wire(0) /=  '0') else MB60_11372;
    -- flow-through select operator MUX_11651_inst
    MC31_11652 <= MB63_11396 when (BITSEL_u8_u1_11648_wire(0) /=  '0') else MB62_11388;
    -- flow-through select operator MUX_11659_inst
    MD0_11660 <= MC1_11412 when (BITSEL_u8_u1_11656_wire(0) /=  '0') else MC0_11404;
    -- flow-through select operator MUX_11667_inst
    MD1_11668 <= MC3_11428 when (BITSEL_u8_u1_11664_wire(0) /=  '0') else MC2_11420;
    -- flow-through select operator MUX_11675_inst
    MD2_11676 <= MC5_11444 when (BITSEL_u8_u1_11672_wire(0) /=  '0') else MC4_11436;
    -- flow-through select operator MUX_11683_inst
    MD3_11684 <= MC7_11460 when (BITSEL_u8_u1_11680_wire(0) /=  '0') else MC6_11452;
    -- flow-through select operator MUX_11691_inst
    MD4_11692 <= MC9_11476 when (BITSEL_u8_u1_11688_wire(0) /=  '0') else MC8_11468;
    -- flow-through select operator MUX_11699_inst
    MD5_11700 <= MC11_11492 when (BITSEL_u8_u1_11696_wire(0) /=  '0') else MC10_11484;
    -- flow-through select operator MUX_11707_inst
    MD6_11708 <= MC13_11508 when (BITSEL_u8_u1_11704_wire(0) /=  '0') else MC12_11500;
    -- flow-through select operator MUX_11715_inst
    MD7_11716 <= MC15_11524 when (BITSEL_u8_u1_11712_wire(0) /=  '0') else MC14_11516;
    -- flow-through select operator MUX_11723_inst
    MD8_11724 <= MC17_11540 when (BITSEL_u8_u1_11720_wire(0) /=  '0') else MC16_11532;
    -- flow-through select operator MUX_11731_inst
    MD9_11732 <= MC19_11556 when (BITSEL_u8_u1_11728_wire(0) /=  '0') else MC18_11548;
    -- flow-through select operator MUX_11739_inst
    MD10_11740 <= MC21_11572 when (BITSEL_u8_u1_11736_wire(0) /=  '0') else MC20_11564;
    -- flow-through select operator MUX_11747_inst
    MD11_11748 <= MC23_11588 when (BITSEL_u8_u1_11744_wire(0) /=  '0') else MC22_11580;
    -- flow-through select operator MUX_11755_inst
    MD12_11756 <= MC25_11604 when (BITSEL_u8_u1_11752_wire(0) /=  '0') else MC24_11596;
    -- flow-through select operator MUX_11763_inst
    MD13_11764 <= MC27_11620 when (BITSEL_u8_u1_11760_wire(0) /=  '0') else MC26_11612;
    -- flow-through select operator MUX_11771_inst
    MD14_11772 <= MC29_11636 when (BITSEL_u8_u1_11768_wire(0) /=  '0') else MC28_11628;
    -- flow-through select operator MUX_11779_inst
    MD15_11780 <= MC31_11652 when (BITSEL_u8_u1_11776_wire(0) /=  '0') else MC30_11644;
    -- flow-through select operator MUX_11787_inst
    ME0_11788 <= MD1_11668 when (BITSEL_u8_u1_11784_wire(0) /=  '0') else MD0_11660;
    -- flow-through select operator MUX_11795_inst
    ME1_11796 <= MD3_11684 when (BITSEL_u8_u1_11792_wire(0) /=  '0') else MD2_11676;
    -- flow-through select operator MUX_11803_inst
    ME2_11804 <= MD5_11700 when (BITSEL_u8_u1_11800_wire(0) /=  '0') else MD4_11692;
    -- flow-through select operator MUX_11811_inst
    ME3_11812 <= MD7_11716 when (BITSEL_u8_u1_11808_wire(0) /=  '0') else MD6_11708;
    -- flow-through select operator MUX_11819_inst
    ME4_11820 <= MD9_11732 when (BITSEL_u8_u1_11816_wire(0) /=  '0') else MD8_11724;
    -- flow-through select operator MUX_11827_inst
    ME5_11828 <= MD11_11748 when (BITSEL_u8_u1_11824_wire(0) /=  '0') else MD10_11740;
    -- flow-through select operator MUX_11835_inst
    ME6_11836 <= MD13_11764 when (BITSEL_u8_u1_11832_wire(0) /=  '0') else MD12_11756;
    -- flow-through select operator MUX_11843_inst
    ME7_11844 <= MD15_11780 when (BITSEL_u8_u1_11840_wire(0) /=  '0') else MD14_11772;
    -- flow-through select operator MUX_11851_inst
    MF0_11852 <= ME1_11796 when (BITSEL_u8_u1_11848_wire(0) /=  '0') else ME0_11788;
    -- flow-through select operator MUX_11859_inst
    MF1_11860 <= ME3_11812 when (BITSEL_u8_u1_11856_wire(0) /=  '0') else ME2_11804;
    -- flow-through select operator MUX_11867_inst
    MF2_11868 <= ME5_11828 when (BITSEL_u8_u1_11864_wire(0) /=  '0') else ME4_11820;
    -- flow-through select operator MUX_11875_inst
    MF3_11876 <= ME7_11844 when (BITSEL_u8_u1_11872_wire(0) /=  '0') else ME6_11836;
    -- flow-through select operator MUX_11883_inst
    MG0_11884 <= MF1_11860 when (BITSEL_u8_u1_11880_wire(0) /=  '0') else MF0_11852;
    -- flow-through select operator MUX_11891_inst
    MG1_11892 <= MF3_11876 when (BITSEL_u8_u1_11888_wire(0) /=  '0') else MF2_11868;
    -- flow-through select operator MUX_11899_inst
    s_out_buffer <= MG1_11892 when (BITSEL_u8_u1_11896_wire(0) /=  '0') else MG0_11884;
    -- flow-through select operator MUX_9613_inst
    MA0_9614 <= type_cast_9610_wire_constant when (BITSEL_u8_u1_9608_wire(0) /=  '0') else type_cast_9612_wire_constant;
    -- flow-through select operator MUX_9623_inst
    MA1_9624 <= type_cast_9620_wire_constant when (BITSEL_u8_u1_9618_wire(0) /=  '0') else type_cast_9622_wire_constant;
    -- flow-through select operator MUX_9633_inst
    MA2_9634 <= type_cast_9630_wire_constant when (BITSEL_u8_u1_9628_wire(0) /=  '0') else type_cast_9632_wire_constant;
    -- flow-through select operator MUX_9643_inst
    MA3_9644 <= type_cast_9640_wire_constant when (BITSEL_u8_u1_9638_wire(0) /=  '0') else type_cast_9642_wire_constant;
    -- flow-through select operator MUX_9653_inst
    MA4_9654 <= type_cast_9650_wire_constant when (BITSEL_u8_u1_9648_wire(0) /=  '0') else type_cast_9652_wire_constant;
    -- flow-through select operator MUX_9663_inst
    MA5_9664 <= type_cast_9660_wire_constant when (BITSEL_u8_u1_9658_wire(0) /=  '0') else type_cast_9662_wire_constant;
    -- flow-through select operator MUX_9673_inst
    MA6_9674 <= type_cast_9670_wire_constant when (BITSEL_u8_u1_9668_wire(0) /=  '0') else type_cast_9672_wire_constant;
    -- flow-through select operator MUX_9683_inst
    MA7_9684 <= type_cast_9680_wire_constant when (BITSEL_u8_u1_9678_wire(0) /=  '0') else type_cast_9682_wire_constant;
    -- flow-through select operator MUX_9693_inst
    MA8_9694 <= type_cast_9690_wire_constant when (BITSEL_u8_u1_9688_wire(0) /=  '0') else type_cast_9692_wire_constant;
    -- flow-through select operator MUX_9703_inst
    MA9_9704 <= type_cast_9700_wire_constant when (BITSEL_u8_u1_9698_wire(0) /=  '0') else type_cast_9702_wire_constant;
    -- flow-through select operator MUX_9713_inst
    MA10_9714 <= type_cast_9710_wire_constant when (BITSEL_u8_u1_9708_wire(0) /=  '0') else type_cast_9712_wire_constant;
    -- flow-through select operator MUX_9723_inst
    MA11_9724 <= type_cast_9720_wire_constant when (BITSEL_u8_u1_9718_wire(0) /=  '0') else type_cast_9722_wire_constant;
    -- flow-through select operator MUX_9733_inst
    MA12_9734 <= type_cast_9730_wire_constant when (BITSEL_u8_u1_9728_wire(0) /=  '0') else type_cast_9732_wire_constant;
    -- flow-through select operator MUX_9743_inst
    MA13_9744 <= type_cast_9740_wire_constant when (BITSEL_u8_u1_9738_wire(0) /=  '0') else type_cast_9742_wire_constant;
    -- flow-through select operator MUX_9753_inst
    MA14_9754 <= type_cast_9750_wire_constant when (BITSEL_u8_u1_9748_wire(0) /=  '0') else type_cast_9752_wire_constant;
    -- flow-through select operator MUX_9763_inst
    MA15_9764 <= type_cast_9760_wire_constant when (BITSEL_u8_u1_9758_wire(0) /=  '0') else type_cast_9762_wire_constant;
    -- flow-through select operator MUX_9773_inst
    MA16_9774 <= type_cast_9770_wire_constant when (BITSEL_u8_u1_9768_wire(0) /=  '0') else type_cast_9772_wire_constant;
    -- flow-through select operator MUX_9783_inst
    MA17_9784 <= type_cast_9780_wire_constant when (BITSEL_u8_u1_9778_wire(0) /=  '0') else type_cast_9782_wire_constant;
    -- flow-through select operator MUX_9793_inst
    MA18_9794 <= type_cast_9790_wire_constant when (BITSEL_u8_u1_9788_wire(0) /=  '0') else type_cast_9792_wire_constant;
    -- flow-through select operator MUX_9803_inst
    MA19_9804 <= type_cast_9800_wire_constant when (BITSEL_u8_u1_9798_wire(0) /=  '0') else type_cast_9802_wire_constant;
    -- flow-through select operator MUX_9813_inst
    MA20_9814 <= type_cast_9810_wire_constant when (BITSEL_u8_u1_9808_wire(0) /=  '0') else type_cast_9812_wire_constant;
    -- flow-through select operator MUX_9823_inst
    MA21_9824 <= type_cast_9820_wire_constant when (BITSEL_u8_u1_9818_wire(0) /=  '0') else type_cast_9822_wire_constant;
    -- flow-through select operator MUX_9833_inst
    MA22_9834 <= type_cast_9830_wire_constant when (BITSEL_u8_u1_9828_wire(0) /=  '0') else type_cast_9832_wire_constant;
    -- flow-through select operator MUX_9843_inst
    MA23_9844 <= type_cast_9840_wire_constant when (BITSEL_u8_u1_9838_wire(0) /=  '0') else type_cast_9842_wire_constant;
    -- flow-through select operator MUX_9853_inst
    MA24_9854 <= type_cast_9850_wire_constant when (BITSEL_u8_u1_9848_wire(0) /=  '0') else type_cast_9852_wire_constant;
    -- flow-through select operator MUX_9863_inst
    MA25_9864 <= type_cast_9860_wire_constant when (BITSEL_u8_u1_9858_wire(0) /=  '0') else type_cast_9862_wire_constant;
    -- flow-through select operator MUX_9873_inst
    MA26_9874 <= type_cast_9870_wire_constant when (BITSEL_u8_u1_9868_wire(0) /=  '0') else type_cast_9872_wire_constant;
    -- flow-through select operator MUX_9883_inst
    MA27_9884 <= type_cast_9880_wire_constant when (BITSEL_u8_u1_9878_wire(0) /=  '0') else type_cast_9882_wire_constant;
    -- flow-through select operator MUX_9893_inst
    MA28_9894 <= type_cast_9890_wire_constant when (BITSEL_u8_u1_9888_wire(0) /=  '0') else type_cast_9892_wire_constant;
    -- flow-through select operator MUX_9903_inst
    MA29_9904 <= type_cast_9900_wire_constant when (BITSEL_u8_u1_9898_wire(0) /=  '0') else type_cast_9902_wire_constant;
    -- flow-through select operator MUX_9913_inst
    MA30_9914 <= type_cast_9910_wire_constant when (BITSEL_u8_u1_9908_wire(0) /=  '0') else type_cast_9912_wire_constant;
    -- flow-through select operator MUX_9923_inst
    MA31_9924 <= type_cast_9920_wire_constant when (BITSEL_u8_u1_9918_wire(0) /=  '0') else type_cast_9922_wire_constant;
    -- flow-through select operator MUX_9933_inst
    MA32_9934 <= type_cast_9930_wire_constant when (BITSEL_u8_u1_9928_wire(0) /=  '0') else type_cast_9932_wire_constant;
    -- flow-through select operator MUX_9943_inst
    MA33_9944 <= type_cast_9940_wire_constant when (BITSEL_u8_u1_9938_wire(0) /=  '0') else type_cast_9942_wire_constant;
    -- flow-through select operator MUX_9953_inst
    MA34_9954 <= type_cast_9950_wire_constant when (BITSEL_u8_u1_9948_wire(0) /=  '0') else type_cast_9952_wire_constant;
    -- flow-through select operator MUX_9963_inst
    MA35_9964 <= type_cast_9960_wire_constant when (BITSEL_u8_u1_9958_wire(0) /=  '0') else type_cast_9962_wire_constant;
    -- flow-through select operator MUX_9973_inst
    MA36_9974 <= type_cast_9970_wire_constant when (BITSEL_u8_u1_9968_wire(0) /=  '0') else type_cast_9972_wire_constant;
    -- flow-through select operator MUX_9983_inst
    MA37_9984 <= type_cast_9980_wire_constant when (BITSEL_u8_u1_9978_wire(0) /=  '0') else type_cast_9982_wire_constant;
    -- flow-through select operator MUX_9993_inst
    MA38_9994 <= type_cast_9990_wire_constant when (BITSEL_u8_u1_9988_wire(0) /=  '0') else type_cast_9992_wire_constant;
    -- binary operator BITSEL_u8_u1_10008_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_10007_wire_constant, tmp_var);
      BITSEL_u8_u1_10008_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_10018_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_10017_wire_constant, tmp_var);
      BITSEL_u8_u1_10018_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_10028_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_10027_wire_constant, tmp_var);
      BITSEL_u8_u1_10028_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_10038_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_10037_wire_constant, tmp_var);
      BITSEL_u8_u1_10038_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_10048_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_10047_wire_constant, tmp_var);
      BITSEL_u8_u1_10048_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_10058_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_10057_wire_constant, tmp_var);
      BITSEL_u8_u1_10058_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_10068_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_10067_wire_constant, tmp_var);
      BITSEL_u8_u1_10068_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_10078_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_10077_wire_constant, tmp_var);
      BITSEL_u8_u1_10078_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_10088_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_10087_wire_constant, tmp_var);
      BITSEL_u8_u1_10088_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_10098_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_10097_wire_constant, tmp_var);
      BITSEL_u8_u1_10098_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_10108_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_10107_wire_constant, tmp_var);
      BITSEL_u8_u1_10108_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_10118_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_10117_wire_constant, tmp_var);
      BITSEL_u8_u1_10118_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_10128_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_10127_wire_constant, tmp_var);
      BITSEL_u8_u1_10128_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_10138_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_10137_wire_constant, tmp_var);
      BITSEL_u8_u1_10138_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_10148_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_10147_wire_constant, tmp_var);
      BITSEL_u8_u1_10148_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_10158_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_10157_wire_constant, tmp_var);
      BITSEL_u8_u1_10158_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_10168_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_10167_wire_constant, tmp_var);
      BITSEL_u8_u1_10168_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_10178_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_10177_wire_constant, tmp_var);
      BITSEL_u8_u1_10178_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_10188_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_10187_wire_constant, tmp_var);
      BITSEL_u8_u1_10188_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_10198_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_10197_wire_constant, tmp_var);
      BITSEL_u8_u1_10198_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_10208_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_10207_wire_constant, tmp_var);
      BITSEL_u8_u1_10208_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_10218_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_10217_wire_constant, tmp_var);
      BITSEL_u8_u1_10218_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_10228_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_10227_wire_constant, tmp_var);
      BITSEL_u8_u1_10228_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_10238_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_10237_wire_constant, tmp_var);
      BITSEL_u8_u1_10238_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_10248_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_10247_wire_constant, tmp_var);
      BITSEL_u8_u1_10248_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_10258_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_10257_wire_constant, tmp_var);
      BITSEL_u8_u1_10258_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_10268_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_10267_wire_constant, tmp_var);
      BITSEL_u8_u1_10268_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_10278_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_10277_wire_constant, tmp_var);
      BITSEL_u8_u1_10278_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_10288_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_10287_wire_constant, tmp_var);
      BITSEL_u8_u1_10288_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_10298_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_10297_wire_constant, tmp_var);
      BITSEL_u8_u1_10298_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_10308_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_10307_wire_constant, tmp_var);
      BITSEL_u8_u1_10308_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_10318_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_10317_wire_constant, tmp_var);
      BITSEL_u8_u1_10318_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_10328_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_10327_wire_constant, tmp_var);
      BITSEL_u8_u1_10328_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_10338_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_10337_wire_constant, tmp_var);
      BITSEL_u8_u1_10338_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_10348_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_10347_wire_constant, tmp_var);
      BITSEL_u8_u1_10348_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_10358_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_10357_wire_constant, tmp_var);
      BITSEL_u8_u1_10358_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_10368_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_10367_wire_constant, tmp_var);
      BITSEL_u8_u1_10368_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_10378_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_10377_wire_constant, tmp_var);
      BITSEL_u8_u1_10378_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_10388_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_10387_wire_constant, tmp_var);
      BITSEL_u8_u1_10388_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_10398_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_10397_wire_constant, tmp_var);
      BITSEL_u8_u1_10398_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_10408_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_10407_wire_constant, tmp_var);
      BITSEL_u8_u1_10408_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_10418_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_10417_wire_constant, tmp_var);
      BITSEL_u8_u1_10418_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_10428_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_10427_wire_constant, tmp_var);
      BITSEL_u8_u1_10428_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_10438_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_10437_wire_constant, tmp_var);
      BITSEL_u8_u1_10438_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_10448_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_10447_wire_constant, tmp_var);
      BITSEL_u8_u1_10448_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_10458_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_10457_wire_constant, tmp_var);
      BITSEL_u8_u1_10458_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_10468_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_10467_wire_constant, tmp_var);
      BITSEL_u8_u1_10468_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_10478_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_10477_wire_constant, tmp_var);
      BITSEL_u8_u1_10478_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_10488_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_10487_wire_constant, tmp_var);
      BITSEL_u8_u1_10488_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_10498_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_10497_wire_constant, tmp_var);
      BITSEL_u8_u1_10498_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_10508_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_10507_wire_constant, tmp_var);
      BITSEL_u8_u1_10508_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_10518_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_10517_wire_constant, tmp_var);
      BITSEL_u8_u1_10518_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_10528_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_10527_wire_constant, tmp_var);
      BITSEL_u8_u1_10528_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_10538_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_10537_wire_constant, tmp_var);
      BITSEL_u8_u1_10538_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_10548_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_10547_wire_constant, tmp_var);
      BITSEL_u8_u1_10548_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_10558_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_10557_wire_constant, tmp_var);
      BITSEL_u8_u1_10558_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_10568_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_10567_wire_constant, tmp_var);
      BITSEL_u8_u1_10568_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_10578_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_10577_wire_constant, tmp_var);
      BITSEL_u8_u1_10578_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_10588_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_10587_wire_constant, tmp_var);
      BITSEL_u8_u1_10588_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_10598_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_10597_wire_constant, tmp_var);
      BITSEL_u8_u1_10598_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_10608_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_10607_wire_constant, tmp_var);
      BITSEL_u8_u1_10608_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_10618_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_10617_wire_constant, tmp_var);
      BITSEL_u8_u1_10618_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_10628_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_10627_wire_constant, tmp_var);
      BITSEL_u8_u1_10628_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_10638_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_10637_wire_constant, tmp_var);
      BITSEL_u8_u1_10638_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_10648_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_10647_wire_constant, tmp_var);
      BITSEL_u8_u1_10648_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_10658_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_10657_wire_constant, tmp_var);
      BITSEL_u8_u1_10658_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_10668_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_10667_wire_constant, tmp_var);
      BITSEL_u8_u1_10668_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_10678_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_10677_wire_constant, tmp_var);
      BITSEL_u8_u1_10678_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_10688_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_10687_wire_constant, tmp_var);
      BITSEL_u8_u1_10688_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_10698_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_10697_wire_constant, tmp_var);
      BITSEL_u8_u1_10698_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_10708_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_10707_wire_constant, tmp_var);
      BITSEL_u8_u1_10708_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_10718_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_10717_wire_constant, tmp_var);
      BITSEL_u8_u1_10718_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_10728_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_10727_wire_constant, tmp_var);
      BITSEL_u8_u1_10728_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_10738_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_10737_wire_constant, tmp_var);
      BITSEL_u8_u1_10738_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_10748_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_10747_wire_constant, tmp_var);
      BITSEL_u8_u1_10748_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_10758_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_10757_wire_constant, tmp_var);
      BITSEL_u8_u1_10758_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_10768_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_10767_wire_constant, tmp_var);
      BITSEL_u8_u1_10768_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_10778_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_10777_wire_constant, tmp_var);
      BITSEL_u8_u1_10778_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_10788_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_10787_wire_constant, tmp_var);
      BITSEL_u8_u1_10788_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_10798_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_10797_wire_constant, tmp_var);
      BITSEL_u8_u1_10798_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_10808_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_10807_wire_constant, tmp_var);
      BITSEL_u8_u1_10808_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_10818_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_10817_wire_constant, tmp_var);
      BITSEL_u8_u1_10818_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_10828_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_10827_wire_constant, tmp_var);
      BITSEL_u8_u1_10828_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_10838_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_10837_wire_constant, tmp_var);
      BITSEL_u8_u1_10838_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_10848_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_10847_wire_constant, tmp_var);
      BITSEL_u8_u1_10848_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_10858_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_10857_wire_constant, tmp_var);
      BITSEL_u8_u1_10858_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_10868_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_10867_wire_constant, tmp_var);
      BITSEL_u8_u1_10868_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_10878_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_10877_wire_constant, tmp_var);
      BITSEL_u8_u1_10878_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_10888_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_10887_wire_constant, tmp_var);
      BITSEL_u8_u1_10888_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_10896_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_10895_wire_constant, tmp_var);
      BITSEL_u8_u1_10896_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_10904_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_10903_wire_constant, tmp_var);
      BITSEL_u8_u1_10904_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_10912_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_10911_wire_constant, tmp_var);
      BITSEL_u8_u1_10912_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_10920_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_10919_wire_constant, tmp_var);
      BITSEL_u8_u1_10920_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_10928_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_10927_wire_constant, tmp_var);
      BITSEL_u8_u1_10928_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_10936_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_10935_wire_constant, tmp_var);
      BITSEL_u8_u1_10936_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_10944_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_10943_wire_constant, tmp_var);
      BITSEL_u8_u1_10944_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_10952_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_10951_wire_constant, tmp_var);
      BITSEL_u8_u1_10952_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_10960_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_10959_wire_constant, tmp_var);
      BITSEL_u8_u1_10960_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_10968_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_10967_wire_constant, tmp_var);
      BITSEL_u8_u1_10968_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_10976_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_10975_wire_constant, tmp_var);
      BITSEL_u8_u1_10976_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_10984_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_10983_wire_constant, tmp_var);
      BITSEL_u8_u1_10984_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_10992_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_10991_wire_constant, tmp_var);
      BITSEL_u8_u1_10992_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11000_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_10999_wire_constant, tmp_var);
      BITSEL_u8_u1_11000_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11008_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11007_wire_constant, tmp_var);
      BITSEL_u8_u1_11008_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11016_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11015_wire_constant, tmp_var);
      BITSEL_u8_u1_11016_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11024_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11023_wire_constant, tmp_var);
      BITSEL_u8_u1_11024_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11032_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11031_wire_constant, tmp_var);
      BITSEL_u8_u1_11032_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11040_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11039_wire_constant, tmp_var);
      BITSEL_u8_u1_11040_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11048_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11047_wire_constant, tmp_var);
      BITSEL_u8_u1_11048_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11056_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11055_wire_constant, tmp_var);
      BITSEL_u8_u1_11056_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11064_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11063_wire_constant, tmp_var);
      BITSEL_u8_u1_11064_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11072_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11071_wire_constant, tmp_var);
      BITSEL_u8_u1_11072_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11080_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11079_wire_constant, tmp_var);
      BITSEL_u8_u1_11080_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11088_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11087_wire_constant, tmp_var);
      BITSEL_u8_u1_11088_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11096_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11095_wire_constant, tmp_var);
      BITSEL_u8_u1_11096_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11104_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11103_wire_constant, tmp_var);
      BITSEL_u8_u1_11104_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11112_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11111_wire_constant, tmp_var);
      BITSEL_u8_u1_11112_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11120_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11119_wire_constant, tmp_var);
      BITSEL_u8_u1_11120_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11128_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11127_wire_constant, tmp_var);
      BITSEL_u8_u1_11128_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11136_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11135_wire_constant, tmp_var);
      BITSEL_u8_u1_11136_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11144_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11143_wire_constant, tmp_var);
      BITSEL_u8_u1_11144_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11152_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11151_wire_constant, tmp_var);
      BITSEL_u8_u1_11152_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11160_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11159_wire_constant, tmp_var);
      BITSEL_u8_u1_11160_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11168_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11167_wire_constant, tmp_var);
      BITSEL_u8_u1_11168_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11176_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11175_wire_constant, tmp_var);
      BITSEL_u8_u1_11176_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11184_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11183_wire_constant, tmp_var);
      BITSEL_u8_u1_11184_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11192_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11191_wire_constant, tmp_var);
      BITSEL_u8_u1_11192_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11200_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11199_wire_constant, tmp_var);
      BITSEL_u8_u1_11200_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11208_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11207_wire_constant, tmp_var);
      BITSEL_u8_u1_11208_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11216_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11215_wire_constant, tmp_var);
      BITSEL_u8_u1_11216_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11224_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11223_wire_constant, tmp_var);
      BITSEL_u8_u1_11224_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11232_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11231_wire_constant, tmp_var);
      BITSEL_u8_u1_11232_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11240_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11239_wire_constant, tmp_var);
      BITSEL_u8_u1_11240_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11248_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11247_wire_constant, tmp_var);
      BITSEL_u8_u1_11248_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11256_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11255_wire_constant, tmp_var);
      BITSEL_u8_u1_11256_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11264_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11263_wire_constant, tmp_var);
      BITSEL_u8_u1_11264_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11272_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11271_wire_constant, tmp_var);
      BITSEL_u8_u1_11272_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11280_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11279_wire_constant, tmp_var);
      BITSEL_u8_u1_11280_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11288_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11287_wire_constant, tmp_var);
      BITSEL_u8_u1_11288_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11296_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11295_wire_constant, tmp_var);
      BITSEL_u8_u1_11296_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11304_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11303_wire_constant, tmp_var);
      BITSEL_u8_u1_11304_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11312_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11311_wire_constant, tmp_var);
      BITSEL_u8_u1_11312_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11320_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11319_wire_constant, tmp_var);
      BITSEL_u8_u1_11320_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11328_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11327_wire_constant, tmp_var);
      BITSEL_u8_u1_11328_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11336_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11335_wire_constant, tmp_var);
      BITSEL_u8_u1_11336_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11344_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11343_wire_constant, tmp_var);
      BITSEL_u8_u1_11344_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11352_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11351_wire_constant, tmp_var);
      BITSEL_u8_u1_11352_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11360_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11359_wire_constant, tmp_var);
      BITSEL_u8_u1_11360_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11368_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11367_wire_constant, tmp_var);
      BITSEL_u8_u1_11368_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11376_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11375_wire_constant, tmp_var);
      BITSEL_u8_u1_11376_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11384_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11383_wire_constant, tmp_var);
      BITSEL_u8_u1_11384_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11392_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11391_wire_constant, tmp_var);
      BITSEL_u8_u1_11392_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11400_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11399_wire_constant, tmp_var);
      BITSEL_u8_u1_11400_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11408_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11407_wire_constant, tmp_var);
      BITSEL_u8_u1_11408_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11416_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11415_wire_constant, tmp_var);
      BITSEL_u8_u1_11416_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11424_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11423_wire_constant, tmp_var);
      BITSEL_u8_u1_11424_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11432_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11431_wire_constant, tmp_var);
      BITSEL_u8_u1_11432_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11440_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11439_wire_constant, tmp_var);
      BITSEL_u8_u1_11440_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11448_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11447_wire_constant, tmp_var);
      BITSEL_u8_u1_11448_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11456_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11455_wire_constant, tmp_var);
      BITSEL_u8_u1_11456_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11464_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11463_wire_constant, tmp_var);
      BITSEL_u8_u1_11464_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11472_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11471_wire_constant, tmp_var);
      BITSEL_u8_u1_11472_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11480_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11479_wire_constant, tmp_var);
      BITSEL_u8_u1_11480_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11488_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11487_wire_constant, tmp_var);
      BITSEL_u8_u1_11488_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11496_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11495_wire_constant, tmp_var);
      BITSEL_u8_u1_11496_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11504_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11503_wire_constant, tmp_var);
      BITSEL_u8_u1_11504_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11512_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11511_wire_constant, tmp_var);
      BITSEL_u8_u1_11512_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11520_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11519_wire_constant, tmp_var);
      BITSEL_u8_u1_11520_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11528_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11527_wire_constant, tmp_var);
      BITSEL_u8_u1_11528_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11536_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11535_wire_constant, tmp_var);
      BITSEL_u8_u1_11536_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11544_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11543_wire_constant, tmp_var);
      BITSEL_u8_u1_11544_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11552_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11551_wire_constant, tmp_var);
      BITSEL_u8_u1_11552_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11560_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11559_wire_constant, tmp_var);
      BITSEL_u8_u1_11560_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11568_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11567_wire_constant, tmp_var);
      BITSEL_u8_u1_11568_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11576_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11575_wire_constant, tmp_var);
      BITSEL_u8_u1_11576_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11584_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11583_wire_constant, tmp_var);
      BITSEL_u8_u1_11584_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11592_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11591_wire_constant, tmp_var);
      BITSEL_u8_u1_11592_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11600_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11599_wire_constant, tmp_var);
      BITSEL_u8_u1_11600_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11608_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11607_wire_constant, tmp_var);
      BITSEL_u8_u1_11608_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11616_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11615_wire_constant, tmp_var);
      BITSEL_u8_u1_11616_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11624_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11623_wire_constant, tmp_var);
      BITSEL_u8_u1_11624_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11632_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11631_wire_constant, tmp_var);
      BITSEL_u8_u1_11632_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11640_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11639_wire_constant, tmp_var);
      BITSEL_u8_u1_11640_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11648_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11647_wire_constant, tmp_var);
      BITSEL_u8_u1_11648_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11656_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11655_wire_constant, tmp_var);
      BITSEL_u8_u1_11656_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11664_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11663_wire_constant, tmp_var);
      BITSEL_u8_u1_11664_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11672_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11671_wire_constant, tmp_var);
      BITSEL_u8_u1_11672_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11680_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11679_wire_constant, tmp_var);
      BITSEL_u8_u1_11680_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11688_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11687_wire_constant, tmp_var);
      BITSEL_u8_u1_11688_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11696_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11695_wire_constant, tmp_var);
      BITSEL_u8_u1_11696_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11704_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11703_wire_constant, tmp_var);
      BITSEL_u8_u1_11704_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11712_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11711_wire_constant, tmp_var);
      BITSEL_u8_u1_11712_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11720_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11719_wire_constant, tmp_var);
      BITSEL_u8_u1_11720_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11728_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11727_wire_constant, tmp_var);
      BITSEL_u8_u1_11728_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11736_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11735_wire_constant, tmp_var);
      BITSEL_u8_u1_11736_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11744_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11743_wire_constant, tmp_var);
      BITSEL_u8_u1_11744_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11752_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11751_wire_constant, tmp_var);
      BITSEL_u8_u1_11752_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11760_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11759_wire_constant, tmp_var);
      BITSEL_u8_u1_11760_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11768_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11767_wire_constant, tmp_var);
      BITSEL_u8_u1_11768_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11776_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11775_wire_constant, tmp_var);
      BITSEL_u8_u1_11776_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11784_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11783_wire_constant, tmp_var);
      BITSEL_u8_u1_11784_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11792_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11791_wire_constant, tmp_var);
      BITSEL_u8_u1_11792_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11800_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11799_wire_constant, tmp_var);
      BITSEL_u8_u1_11800_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11808_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11807_wire_constant, tmp_var);
      BITSEL_u8_u1_11808_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11816_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11815_wire_constant, tmp_var);
      BITSEL_u8_u1_11816_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11824_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11823_wire_constant, tmp_var);
      BITSEL_u8_u1_11824_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11832_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11831_wire_constant, tmp_var);
      BITSEL_u8_u1_11832_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11840_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11839_wire_constant, tmp_var);
      BITSEL_u8_u1_11840_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11848_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11847_wire_constant, tmp_var);
      BITSEL_u8_u1_11848_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11856_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11855_wire_constant, tmp_var);
      BITSEL_u8_u1_11856_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11864_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11863_wire_constant, tmp_var);
      BITSEL_u8_u1_11864_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11872_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11871_wire_constant, tmp_var);
      BITSEL_u8_u1_11872_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11880_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11879_wire_constant, tmp_var);
      BITSEL_u8_u1_11880_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11888_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11887_wire_constant, tmp_var);
      BITSEL_u8_u1_11888_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_11896_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_11895_wire_constant, tmp_var);
      BITSEL_u8_u1_11896_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_9608_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_9607_wire_constant, tmp_var);
      BITSEL_u8_u1_9608_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_9618_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_9617_wire_constant, tmp_var);
      BITSEL_u8_u1_9618_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_9628_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_9627_wire_constant, tmp_var);
      BITSEL_u8_u1_9628_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_9638_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_9637_wire_constant, tmp_var);
      BITSEL_u8_u1_9638_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_9648_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_9647_wire_constant, tmp_var);
      BITSEL_u8_u1_9648_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_9658_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_9657_wire_constant, tmp_var);
      BITSEL_u8_u1_9658_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_9668_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_9667_wire_constant, tmp_var);
      BITSEL_u8_u1_9668_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_9678_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_9677_wire_constant, tmp_var);
      BITSEL_u8_u1_9678_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_9688_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_9687_wire_constant, tmp_var);
      BITSEL_u8_u1_9688_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_9698_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_9697_wire_constant, tmp_var);
      BITSEL_u8_u1_9698_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_9708_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_9707_wire_constant, tmp_var);
      BITSEL_u8_u1_9708_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_9718_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_9717_wire_constant, tmp_var);
      BITSEL_u8_u1_9718_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_9728_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_9727_wire_constant, tmp_var);
      BITSEL_u8_u1_9728_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_9738_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_9737_wire_constant, tmp_var);
      BITSEL_u8_u1_9738_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_9748_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_9747_wire_constant, tmp_var);
      BITSEL_u8_u1_9748_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_9758_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_9757_wire_constant, tmp_var);
      BITSEL_u8_u1_9758_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_9768_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_9767_wire_constant, tmp_var);
      BITSEL_u8_u1_9768_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_9778_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_9777_wire_constant, tmp_var);
      BITSEL_u8_u1_9778_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_9788_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_9787_wire_constant, tmp_var);
      BITSEL_u8_u1_9788_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_9798_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_9797_wire_constant, tmp_var);
      BITSEL_u8_u1_9798_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_9808_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_9807_wire_constant, tmp_var);
      BITSEL_u8_u1_9808_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_9818_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_9817_wire_constant, tmp_var);
      BITSEL_u8_u1_9818_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_9828_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_9827_wire_constant, tmp_var);
      BITSEL_u8_u1_9828_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_9838_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_9837_wire_constant, tmp_var);
      BITSEL_u8_u1_9838_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_9848_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_9847_wire_constant, tmp_var);
      BITSEL_u8_u1_9848_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_9858_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_9857_wire_constant, tmp_var);
      BITSEL_u8_u1_9858_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_9868_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_9867_wire_constant, tmp_var);
      BITSEL_u8_u1_9868_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_9878_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_9877_wire_constant, tmp_var);
      BITSEL_u8_u1_9878_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_9888_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_9887_wire_constant, tmp_var);
      BITSEL_u8_u1_9888_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_9898_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_9897_wire_constant, tmp_var);
      BITSEL_u8_u1_9898_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_9908_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_9907_wire_constant, tmp_var);
      BITSEL_u8_u1_9908_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_9918_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_9917_wire_constant, tmp_var);
      BITSEL_u8_u1_9918_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_9928_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_9927_wire_constant, tmp_var);
      BITSEL_u8_u1_9928_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_9938_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_9937_wire_constant, tmp_var);
      BITSEL_u8_u1_9938_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_9948_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_9947_wire_constant, tmp_var);
      BITSEL_u8_u1_9948_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_9958_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_9957_wire_constant, tmp_var);
      BITSEL_u8_u1_9958_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_9968_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_9967_wire_constant, tmp_var);
      BITSEL_u8_u1_9968_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_9978_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_9977_wire_constant, tmp_var);
      BITSEL_u8_u1_9978_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_9988_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_9987_wire_constant, tmp_var);
      BITSEL_u8_u1_9988_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_9998_inst
    process(data_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(data_in_buffer, konst_9997_wire_constant, tmp_var);
      BITSEL_u8_u1_9998_wire <= tmp_var; -- 
    end process;
    -- 
  end Block; -- data_path
  -- 
end sbox_mux_impl_Volatile_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library work;
use work.ahir_system_global_package.all;
entity w_in_buff_daemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    in_data_pipe_read_req : out  std_logic_vector(0 downto 0);
    in_data_pipe_read_ack : in   std_logic_vector(0 downto 0);
    in_data_pipe_read_data : in   std_logic_vector(63 downto 0);
    w_in_buf_pipe_write_req : out  std_logic_vector(0 downto 0);
    w_in_buf_pipe_write_ack : in   std_logic_vector(0 downto 0);
    w_in_buf_pipe_write_data : out  std_logic_vector(127 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity w_in_buff_daemon;
architecture w_in_buff_daemon_arch of w_in_buff_daemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal w_in_buff_daemon_CP_12370_start: Boolean;
  signal w_in_buff_daemon_CP_12370_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal RPIPE_in_data_13974_inst_req_0 : boolean;
  signal RPIPE_in_data_13974_inst_ack_0 : boolean;
  signal RPIPE_in_data_13977_inst_ack_0 : boolean;
  signal do_while_stmt_13971_branch_req_0 : boolean;
  signal RPIPE_in_data_13977_inst_req_0 : boolean;
  signal RPIPE_in_data_13974_inst_ack_1 : boolean;
  signal RPIPE_in_data_13974_inst_req_1 : boolean;
  signal RPIPE_in_data_13977_inst_ack_1 : boolean;
  signal RPIPE_in_data_13977_inst_req_1 : boolean;
  signal do_while_stmt_13971_branch_ack_1 : boolean;
  signal do_while_stmt_13971_branch_ack_0 : boolean;
  signal WPIPE_w_in_buf_13979_inst_ack_1 : boolean;
  signal WPIPE_w_in_buf_13979_inst_req_1 : boolean;
  signal WPIPE_w_in_buf_13979_inst_ack_0 : boolean;
  signal WPIPE_w_in_buf_13979_inst_req_0 : boolean;
  signal CONCAT_u64_u128_13982_inst_ack_1 : boolean;
  signal CONCAT_u64_u128_13982_inst_req_1 : boolean;
  signal CONCAT_u64_u128_13982_inst_ack_0 : boolean;
  signal CONCAT_u64_u128_13982_inst_req_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "w_in_buff_daemon_input_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      bypass_flag => true,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  w_in_buff_daemon_CP_12370_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "w_in_buff_daemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= w_in_buff_daemon_CP_12370_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= w_in_buff_daemon_CP_12370_start & tag_ilock_write_ack_symbol;
    gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= w_in_buff_daemon_CP_12370_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  w_in_buff_daemon_CP_12370: Block -- control-path 
    signal w_in_buff_daemon_CP_12370_elements: BooleanArray(33 downto 0);
    -- 
  begin -- 
    w_in_buff_daemon_CP_12370_elements(0) <= w_in_buff_daemon_CP_12370_start;
    w_in_buff_daemon_CP_12370_symbol <= w_in_buff_daemon_CP_12370_elements(33);
    -- CP-element group 0:  transition  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (2) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_13970/$entry
      -- 
    -- CP-element group 1:  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	3 
    -- CP-element group 1:  members (2) 
      -- CP-element group 1: 	 branch_block_stmt_13970/branch_block_stmt_13970__entry__
      -- CP-element group 1: 	 branch_block_stmt_13970/do_while_stmt_13971__entry__
      -- 
    w_in_buff_daemon_CP_12370_elements(1) <= w_in_buff_daemon_CP_12370_elements(0);
    -- CP-element group 2:  place  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	32 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	33 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_13970/branch_block_stmt_13970__exit__
      -- CP-element group 2: 	 branch_block_stmt_13970/do_while_stmt_13971__exit__
      -- 
    w_in_buff_daemon_CP_12370_elements(2) <= w_in_buff_daemon_CP_12370_elements(32);
    -- CP-element group 3:  transition  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	1 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_13970/do_while_stmt_13971/$entry
      -- 
    w_in_buff_daemon_CP_12370_elements(3) <= w_in_buff_daemon_CP_12370_elements(1);
    -- CP-element group 4:  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	10 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_13970/do_while_stmt_13971/do_while_stmt_13971__entry__
      -- 
    w_in_buff_daemon_CP_12370_elements(4) <= w_in_buff_daemon_CP_12370_elements(3);
    -- CP-element group 5:  merge  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	32 
    -- CP-element group 5:  members (1) 
      -- CP-element group 5: 	 branch_block_stmt_13970/do_while_stmt_13971/do_while_stmt_13971__exit__
      -- 
    -- Element group w_in_buff_daemon_CP_12370_elements(5) is bound as output of CP function.
    -- CP-element group 6:  merge  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	9 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_13970/do_while_stmt_13971/loop_back
      -- 
    -- Element group w_in_buff_daemon_CP_12370_elements(6) is bound as output of CP function.
    -- CP-element group 7:  branch  place  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	11 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	30 
    -- CP-element group 7: 	28 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_13970/do_while_stmt_13971/condition_done
      -- 
    w_in_buff_daemon_CP_12370_elements(7) <= w_in_buff_daemon_CP_12370_elements(11);
    -- CP-element group 8:  branch  place  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	27 
    -- CP-element group 8: successors 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_13970/do_while_stmt_13971/loop_body_done
      -- 
    w_in_buff_daemon_CP_12370_elements(8) <= w_in_buff_daemon_CP_12370_elements(27);
    -- CP-element group 9:  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	6 
    -- CP-element group 9: successors 
    -- CP-element group 9:  members (1) 
      -- CP-element group 9: 	 branch_block_stmt_13970/do_while_stmt_13971/do_while_stmt_13971_loop_body/back_edge_to_loop_body
      -- 
    w_in_buff_daemon_CP_12370_elements(9) <= w_in_buff_daemon_CP_12370_elements(6);
    -- CP-element group 10:  transition  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	4 
    -- CP-element group 10: successors 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_13970/do_while_stmt_13971/do_while_stmt_13971_loop_body/first_time_through_loop_body
      -- 
    w_in_buff_daemon_CP_12370_elements(10) <= w_in_buff_daemon_CP_12370_elements(4);
    -- CP-element group 11:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	21 
    -- CP-element group 11: 	7 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 branch_block_stmt_13970/do_while_stmt_13971/do_while_stmt_13971_loop_body/$entry
      -- CP-element group 11: 	 branch_block_stmt_13970/do_while_stmt_13971/do_while_stmt_13971_loop_body/loop_body_start
      -- CP-element group 11: 	 branch_block_stmt_13970/do_while_stmt_13971/do_while_stmt_13971_loop_body/condition_evaluated
      -- 
    condition_evaluated_12394_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_12394_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => w_in_buff_daemon_CP_12370_elements(11), ack => do_while_stmt_13971_branch_req_0); -- 
    -- Element group w_in_buff_daemon_CP_12370_elements(11) is bound as output of CP function.
    -- CP-element group 12:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: marked-predecessors 
    -- CP-element group 12: 	14 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	14 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_13970/do_while_stmt_13971/do_while_stmt_13971_loop_body/RPIPE_in_data_13974_Sample/rr
      -- CP-element group 12: 	 branch_block_stmt_13970/do_while_stmt_13971/do_while_stmt_13971_loop_body/RPIPE_in_data_13974_sample_start_
      -- CP-element group 12: 	 branch_block_stmt_13970/do_while_stmt_13971/do_while_stmt_13971_loop_body/RPIPE_in_data_13974_Sample/$entry
      -- 
    rr_12403_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_12403_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => w_in_buff_daemon_CP_12370_elements(12), ack => RPIPE_in_data_13974_inst_req_0); -- 
    w_in_buff_daemon_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 36) := "w_in_buff_daemon_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= w_in_buff_daemon_CP_12370_elements(11) & w_in_buff_daemon_CP_12370_elements(14);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => w_in_buff_daemon_CP_12370_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	14 
    -- CP-element group 13: marked-predecessors 
    -- CP-element group 13: 	22 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	15 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 branch_block_stmt_13970/do_while_stmt_13971/do_while_stmt_13971_loop_body/RPIPE_in_data_13974_Update/$entry
      -- CP-element group 13: 	 branch_block_stmt_13970/do_while_stmt_13971/do_while_stmt_13971_loop_body/RPIPE_in_data_13974_Update/cr
      -- CP-element group 13: 	 branch_block_stmt_13970/do_while_stmt_13971/do_while_stmt_13971_loop_body/RPIPE_in_data_13974_update_start_
      -- 
    cr_12408_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_12408_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => w_in_buff_daemon_CP_12370_elements(13), ack => RPIPE_in_data_13974_inst_req_1); -- 
    w_in_buff_daemon_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 36) := "w_in_buff_daemon_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= w_in_buff_daemon_CP_12370_elements(14) & w_in_buff_daemon_CP_12370_elements(22);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => w_in_buff_daemon_CP_12370_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	12 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	12 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_13970/do_while_stmt_13971/do_while_stmt_13971_loop_body/RPIPE_in_data_13974_Sample/$exit
      -- CP-element group 14: 	 branch_block_stmt_13970/do_while_stmt_13971/do_while_stmt_13971_loop_body/RPIPE_in_data_13974_Sample/ra
      -- CP-element group 14: 	 branch_block_stmt_13970/do_while_stmt_13971/do_while_stmt_13971_loop_body/RPIPE_in_data_13974_sample_completed_
      -- 
    ra_12404_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_in_data_13974_inst_ack_0, ack => w_in_buff_daemon_CP_12370_elements(14)); -- 
    -- CP-element group 15:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	13 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15: 	20 
    -- CP-element group 15:  members (7) 
      -- CP-element group 15: 	 branch_block_stmt_13970/do_while_stmt_13971/do_while_stmt_13971_loop_body/R_Ina_13980_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_13970/do_while_stmt_13971/do_while_stmt_13971_loop_body/R_Ina_13980_update_start_
      -- CP-element group 15: 	 branch_block_stmt_13970/do_while_stmt_13971/do_while_stmt_13971_loop_body/RPIPE_in_data_13974_Update/ca
      -- CP-element group 15: 	 branch_block_stmt_13970/do_while_stmt_13971/do_while_stmt_13971_loop_body/RPIPE_in_data_13974_Update/$exit
      -- CP-element group 15: 	 branch_block_stmt_13970/do_while_stmt_13971/do_while_stmt_13971_loop_body/RPIPE_in_data_13974_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_13970/do_while_stmt_13971/do_while_stmt_13971_loop_body/R_Ina_13980_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_13970/do_while_stmt_13971/do_while_stmt_13971_loop_body/R_Ina_13980_update_completed_
      -- 
    ca_12409_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_in_data_13974_inst_ack_1, ack => w_in_buff_daemon_CP_12370_elements(15)); -- 
    -- CP-element group 16:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	18 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	18 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_13970/do_while_stmt_13971/do_while_stmt_13971_loop_body/RPIPE_in_data_13977_Sample/rr
      -- CP-element group 16: 	 branch_block_stmt_13970/do_while_stmt_13971/do_while_stmt_13971_loop_body/RPIPE_in_data_13977_Sample/$entry
      -- CP-element group 16: 	 branch_block_stmt_13970/do_while_stmt_13971/do_while_stmt_13971_loop_body/RPIPE_in_data_13977_sample_start_
      -- 
    rr_12417_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_12417_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => w_in_buff_daemon_CP_12370_elements(16), ack => RPIPE_in_data_13977_inst_req_0); -- 
    w_in_buff_daemon_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 36) := "w_in_buff_daemon_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= w_in_buff_daemon_CP_12370_elements(15) & w_in_buff_daemon_CP_12370_elements(18);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => w_in_buff_daemon_CP_12370_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	18 
    -- CP-element group 17: marked-predecessors 
    -- CP-element group 17: 	22 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	19 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 branch_block_stmt_13970/do_while_stmt_13971/do_while_stmt_13971_loop_body/RPIPE_in_data_13977_update_start_
      -- CP-element group 17: 	 branch_block_stmt_13970/do_while_stmt_13971/do_while_stmt_13971_loop_body/RPIPE_in_data_13977_Update/$entry
      -- CP-element group 17: 	 branch_block_stmt_13970/do_while_stmt_13971/do_while_stmt_13971_loop_body/RPIPE_in_data_13977_Update/cr
      -- 
    cr_12422_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_12422_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => w_in_buff_daemon_CP_12370_elements(17), ack => RPIPE_in_data_13977_inst_req_1); -- 
    w_in_buff_daemon_cp_element_group_17: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 36) := "w_in_buff_daemon_cp_element_group_17"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= w_in_buff_daemon_CP_12370_elements(18) & w_in_buff_daemon_CP_12370_elements(22);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => w_in_buff_daemon_CP_12370_elements(17), clk => clk, reset => reset); --
    end block;
    -- CP-element group 18:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	16 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: marked-successors 
    -- CP-element group 18: 	16 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 branch_block_stmt_13970/do_while_stmt_13971/do_while_stmt_13971_loop_body/RPIPE_in_data_13977_sample_completed_
      -- CP-element group 18: 	 branch_block_stmt_13970/do_while_stmt_13971/do_while_stmt_13971_loop_body/RPIPE_in_data_13977_Sample/ra
      -- CP-element group 18: 	 branch_block_stmt_13970/do_while_stmt_13971/do_while_stmt_13971_loop_body/RPIPE_in_data_13977_Sample/$exit
      -- 
    ra_12418_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_in_data_13977_inst_ack_0, ack => w_in_buff_daemon_CP_12370_elements(18)); -- 
    -- CP-element group 19:  transition  input  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	17 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19:  members (7) 
      -- CP-element group 19: 	 branch_block_stmt_13970/do_while_stmt_13971/do_while_stmt_13971_loop_body/RPIPE_in_data_13977_update_completed_
      -- CP-element group 19: 	 branch_block_stmt_13970/do_while_stmt_13971/do_while_stmt_13971_loop_body/RPIPE_in_data_13977_Update/ca
      -- CP-element group 19: 	 branch_block_stmt_13970/do_while_stmt_13971/do_while_stmt_13971_loop_body/RPIPE_in_data_13977_Update/$exit
      -- CP-element group 19: 	 branch_block_stmt_13970/do_while_stmt_13971/do_while_stmt_13971_loop_body/R_Inb_13981_update_completed_
      -- CP-element group 19: 	 branch_block_stmt_13970/do_while_stmt_13971/do_while_stmt_13971_loop_body/R_Inb_13981_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_13970/do_while_stmt_13971/do_while_stmt_13971_loop_body/R_Inb_13981_update_start_
      -- CP-element group 19: 	 branch_block_stmt_13970/do_while_stmt_13971/do_while_stmt_13971_loop_body/R_Inb_13981_sample_start_
      -- 
    ca_12423_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_in_data_13977_inst_ack_1, ack => w_in_buff_daemon_CP_12370_elements(19)); -- 
    -- CP-element group 20:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	15 
    -- CP-element group 20: 	19 
    -- CP-element group 20: marked-predecessors 
    -- CP-element group 20: 	22 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	22 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_13970/do_while_stmt_13971/do_while_stmt_13971_loop_body/CONCAT_u64_u128_13982_sample_start_
      -- CP-element group 20: 	 branch_block_stmt_13970/do_while_stmt_13971/do_while_stmt_13971_loop_body/CONCAT_u64_u128_13982_Sample/rr
      -- CP-element group 20: 	 branch_block_stmt_13970/do_while_stmt_13971/do_while_stmt_13971_loop_body/CONCAT_u64_u128_13982_Sample/$entry
      -- 
    rr_12439_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_12439_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => w_in_buff_daemon_CP_12370_elements(20), ack => CONCAT_u64_u128_13982_inst_req_0); -- 
    w_in_buff_daemon_cp_element_group_20: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 3,1 => 3,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 36) := "w_in_buff_daemon_cp_element_group_20"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= w_in_buff_daemon_CP_12370_elements(15) & w_in_buff_daemon_CP_12370_elements(19) & w_in_buff_daemon_CP_12370_elements(22);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => w_in_buff_daemon_CP_12370_elements(20), clk => clk, reset => reset); --
    end block;
    -- CP-element group 21:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	11 
    -- CP-element group 21: marked-predecessors 
    -- CP-element group 21: 	26 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	23 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_13970/do_while_stmt_13971/do_while_stmt_13971_loop_body/CONCAT_u64_u128_13982_update_start_
      -- CP-element group 21: 	 branch_block_stmt_13970/do_while_stmt_13971/do_while_stmt_13971_loop_body/CONCAT_u64_u128_13982_Update/$entry
      -- CP-element group 21: 	 branch_block_stmt_13970/do_while_stmt_13971/do_while_stmt_13971_loop_body/CONCAT_u64_u128_13982_Update/cr
      -- 
    cr_12444_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_12444_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => w_in_buff_daemon_CP_12370_elements(21), ack => CONCAT_u64_u128_13982_inst_req_1); -- 
    w_in_buff_daemon_cp_element_group_21: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 36) := "w_in_buff_daemon_cp_element_group_21"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= w_in_buff_daemon_CP_12370_elements(11) & w_in_buff_daemon_CP_12370_elements(26);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => w_in_buff_daemon_CP_12370_elements(21), clk => clk, reset => reset); --
    end block;
    -- CP-element group 22:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	20 
    -- CP-element group 22: successors 
    -- CP-element group 22: marked-successors 
    -- CP-element group 22: 	13 
    -- CP-element group 22: 	17 
    -- CP-element group 22: 	20 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_13970/do_while_stmt_13971/do_while_stmt_13971_loop_body/CONCAT_u64_u128_13982_sample_completed_
      -- CP-element group 22: 	 branch_block_stmt_13970/do_while_stmt_13971/do_while_stmt_13971_loop_body/CONCAT_u64_u128_13982_Sample/ra
      -- CP-element group 22: 	 branch_block_stmt_13970/do_while_stmt_13971/do_while_stmt_13971_loop_body/CONCAT_u64_u128_13982_Sample/$exit
      -- 
    ra_12440_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u64_u128_13982_inst_ack_0, ack => w_in_buff_daemon_CP_12370_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	21 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	24 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_13970/do_while_stmt_13971/do_while_stmt_13971_loop_body/CONCAT_u64_u128_13982_update_completed_
      -- CP-element group 23: 	 branch_block_stmt_13970/do_while_stmt_13971/do_while_stmt_13971_loop_body/CONCAT_u64_u128_13982_Update/ca
      -- CP-element group 23: 	 branch_block_stmt_13970/do_while_stmt_13971/do_while_stmt_13971_loop_body/CONCAT_u64_u128_13982_Update/$exit
      -- 
    ca_12445_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u64_u128_13982_inst_ack_1, ack => w_in_buff_daemon_CP_12370_elements(23)); -- 
    -- CP-element group 24:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	23 
    -- CP-element group 24: marked-predecessors 
    -- CP-element group 24: 	26 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	26 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_13970/do_while_stmt_13971/do_while_stmt_13971_loop_body/WPIPE_w_in_buf_13979_Sample/$entry
      -- CP-element group 24: 	 branch_block_stmt_13970/do_while_stmt_13971/do_while_stmt_13971_loop_body/WPIPE_w_in_buf_13979_Sample/req
      -- CP-element group 24: 	 branch_block_stmt_13970/do_while_stmt_13971/do_while_stmt_13971_loop_body/WPIPE_w_in_buf_13979_sample_start_
      -- 
    req_12453_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_12453_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => w_in_buff_daemon_CP_12370_elements(24), ack => WPIPE_w_in_buf_13979_inst_req_0); -- 
    w_in_buff_daemon_cp_element_group_24: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 36) := "w_in_buff_daemon_cp_element_group_24"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= w_in_buff_daemon_CP_12370_elements(23) & w_in_buff_daemon_CP_12370_elements(26);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => w_in_buff_daemon_CP_12370_elements(24), clk => clk, reset => reset); --
    end block;
    -- CP-element group 25:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	26 
    -- CP-element group 25: marked-predecessors 
    -- CP-element group 25: 	27 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	27 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 branch_block_stmt_13970/do_while_stmt_13971/do_while_stmt_13971_loop_body/WPIPE_w_in_buf_13979_Update/$entry
      -- CP-element group 25: 	 branch_block_stmt_13970/do_while_stmt_13971/do_while_stmt_13971_loop_body/WPIPE_w_in_buf_13979_Update/req
      -- CP-element group 25: 	 branch_block_stmt_13970/do_while_stmt_13971/do_while_stmt_13971_loop_body/WPIPE_w_in_buf_13979_update_start_
      -- 
    req_12458_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_12458_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => w_in_buff_daemon_CP_12370_elements(25), ack => WPIPE_w_in_buf_13979_inst_req_1); -- 
    w_in_buff_daemon_cp_element_group_25: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 36) := "w_in_buff_daemon_cp_element_group_25"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= w_in_buff_daemon_CP_12370_elements(26) & w_in_buff_daemon_CP_12370_elements(27);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => w_in_buff_daemon_CP_12370_elements(25), clk => clk, reset => reset); --
    end block;
    -- CP-element group 26:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	24 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	25 
    -- CP-element group 26: marked-successors 
    -- CP-element group 26: 	21 
    -- CP-element group 26: 	24 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_13970/do_while_stmt_13971/do_while_stmt_13971_loop_body/WPIPE_w_in_buf_13979_Sample/ack
      -- CP-element group 26: 	 branch_block_stmt_13970/do_while_stmt_13971/do_while_stmt_13971_loop_body/WPIPE_w_in_buf_13979_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_13970/do_while_stmt_13971/do_while_stmt_13971_loop_body/WPIPE_w_in_buf_13979_sample_completed_
      -- 
    ack_12454_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_w_in_buf_13979_inst_ack_0, ack => w_in_buff_daemon_CP_12370_elements(26)); -- 
    -- CP-element group 27:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	25 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	8 
    -- CP-element group 27: marked-successors 
    -- CP-element group 27: 	25 
    -- CP-element group 27:  members (4) 
      -- CP-element group 27: 	 branch_block_stmt_13970/do_while_stmt_13971/do_while_stmt_13971_loop_body/$exit
      -- CP-element group 27: 	 branch_block_stmt_13970/do_while_stmt_13971/do_while_stmt_13971_loop_body/WPIPE_w_in_buf_13979_Update/ack
      -- CP-element group 27: 	 branch_block_stmt_13970/do_while_stmt_13971/do_while_stmt_13971_loop_body/WPIPE_w_in_buf_13979_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_13970/do_while_stmt_13971/do_while_stmt_13971_loop_body/WPIPE_w_in_buf_13979_update_completed_
      -- 
    ack_12459_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_w_in_buf_13979_inst_ack_1, ack => w_in_buff_daemon_CP_12370_elements(27)); -- 
    -- CP-element group 28:  transition  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	7 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28:  members (1) 
      -- CP-element group 28: 	 branch_block_stmt_13970/do_while_stmt_13971/loop_exit/$entry
      -- 
    w_in_buff_daemon_CP_12370_elements(28) <= w_in_buff_daemon_CP_12370_elements(7);
    -- CP-element group 29:  transition  input  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	28 
    -- CP-element group 29: successors 
    -- CP-element group 29:  members (2) 
      -- CP-element group 29: 	 branch_block_stmt_13970/do_while_stmt_13971/loop_exit/$exit
      -- CP-element group 29: 	 branch_block_stmt_13970/do_while_stmt_13971/loop_exit/ack
      -- 
    ack_12463_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_13971_branch_ack_0, ack => w_in_buff_daemon_CP_12370_elements(29)); -- 
    -- CP-element group 30:  transition  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	7 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30:  members (1) 
      -- CP-element group 30: 	 branch_block_stmt_13970/do_while_stmt_13971/loop_taken/$entry
      -- 
    w_in_buff_daemon_CP_12370_elements(30) <= w_in_buff_daemon_CP_12370_elements(7);
    -- CP-element group 31:  transition  input  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (2) 
      -- CP-element group 31: 	 branch_block_stmt_13970/do_while_stmt_13971/loop_taken/$exit
      -- CP-element group 31: 	 branch_block_stmt_13970/do_while_stmt_13971/loop_taken/ack
      -- 
    ack_12467_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_13971_branch_ack_1, ack => w_in_buff_daemon_CP_12370_elements(31)); -- 
    -- CP-element group 32:  transition  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	5 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	2 
    -- CP-element group 32:  members (1) 
      -- CP-element group 32: 	 branch_block_stmt_13970/do_while_stmt_13971/$exit
      -- 
    w_in_buff_daemon_CP_12370_elements(32) <= w_in_buff_daemon_CP_12370_elements(5);
    -- CP-element group 33:  transition  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	2 
    -- CP-element group 33: successors 
    -- CP-element group 33:  members (2) 
      -- CP-element group 33: 	 $exit
      -- CP-element group 33: 	 branch_block_stmt_13970/$exit
      -- 
    w_in_buff_daemon_CP_12370_elements(33) <= w_in_buff_daemon_CP_12370_elements(2);
    do_while_stmt_13971_terminator_12468: loop_terminator -- 
      generic map (name => " do_while_stmt_13971_terminator_12468", max_iterations_in_flight =>3) 
      port map(loop_body_exit => w_in_buff_daemon_CP_12370_elements(8),loop_continue => w_in_buff_daemon_CP_12370_elements(31),loop_terminate => w_in_buff_daemon_CP_12370_elements(29),loop_back => w_in_buff_daemon_CP_12370_elements(6),loop_exit => w_in_buff_daemon_CP_12370_elements(5),clk => clk, reset => reset); -- 
    entry_tmerge_12395_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= w_in_buff_daemon_CP_12370_elements(9);
        preds(1)  <= w_in_buff_daemon_CP_12370_elements(10);
        entry_tmerge_12395 : transition_merge -- 
          generic map(name => " entry_tmerge_12395")
          port map (preds => preds, symbol_out => w_in_buff_daemon_CP_12370_elements(11));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal CONCAT_u64_u128_13982_wire : std_logic_vector(127 downto 0);
    signal Ina_13975 : std_logic_vector(63 downto 0);
    signal Inb_13978 : std_logic_vector(63 downto 0);
    signal konst_13985_wire_constant : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    konst_13985_wire_constant <= "1";
    do_while_stmt_13971_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= konst_13985_wire_constant;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_13971_branch", condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_13971_branch_req_0,
          ack0 => do_while_stmt_13971_branch_ack_0,
          ack1 => do_while_stmt_13971_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- shared split operator group (0) : CONCAT_u64_u128_13982_inst 
    ApConcat_group_0: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= Ina_13975 & Inb_13978;
      CONCAT_u64_u128_13982_wire <= data_out(127 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= CONCAT_u64_u128_13982_inst_req_0;
      CONCAT_u64_u128_13982_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= CONCAT_u64_u128_13982_inst_req_1;
      CONCAT_u64_u128_13982_inst_ack_1 <= ackR_unguarded(0);
      gI: SplitGuardInterface generic map(name => "gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApConcat",
          name => "ApConcat_group_0",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 64, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 128,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- shared inport operator group (0) : RPIPE_in_data_13977_inst RPIPE_in_data_13974_inst 
    InportGroup0: Block -- 
      signal data_out: std_logic_vector(127 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 1 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 2, 0 => 2);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= RPIPE_in_data_13977_inst_req_0;
      reqL_unguarded(0) <= RPIPE_in_data_13974_inst_req_0;
      RPIPE_in_data_13977_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_in_data_13974_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= RPIPE_in_data_13977_inst_req_1;
      reqR_unguarded(0) <= RPIPE_in_data_13974_inst_req_1;
      RPIPE_in_data_13977_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_in_data_13974_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      gI: SplitGuardInterface generic map(name => "gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Inb_13978 <= data_out(127 downto 64);
      Ina_13975 <= data_out(63 downto 0);
      in_data_read_0: InputPortRevised -- 
        generic map ( name => "in_data_read_0", data_width => 64,  num_reqs => 2,  output_buffering => outBUFs,   no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => in_data_pipe_read_req(0),
          oack => in_data_pipe_read_ack(0),
          odata => in_data_pipe_read_data(63 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_w_in_buf_13979_inst 
    OutportGroup0: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_w_in_buf_13979_inst_req_0;
      WPIPE_w_in_buf_13979_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_w_in_buf_13979_inst_req_1;
      WPIPE_w_in_buf_13979_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      gI: SplitGuardInterface generic map(name => "gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      data_in <= CONCAT_u64_u128_13982_wire;
      w_in_buf_write_0: OutputPortRevised -- 
        generic map ( name => "w_in_buf", data_width => 128, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => w_in_buf_pipe_write_req(0),
          oack => w_in_buf_pipe_write_ack(0),
          odata => w_in_buf_pipe_write_data(127 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end w_in_buff_daemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library work;
use work.ahir_system_global_package.all;
entity w_out_buff_daemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    w_out_buf_pipe_read_req : out  std_logic_vector(0 downto 0);
    w_out_buf_pipe_read_ack : in   std_logic_vector(0 downto 0);
    w_out_buf_pipe_read_data : in   std_logic_vector(127 downto 0);
    out_data_pipe_write_req : out  std_logic_vector(0 downto 0);
    out_data_pipe_write_ack : in   std_logic_vector(0 downto 0);
    out_data_pipe_write_data : out  std_logic_vector(63 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity w_out_buff_daemon;
architecture w_out_buff_daemon_arch of w_out_buff_daemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal w_out_buff_daemon_CP_12469_start: Boolean;
  signal w_out_buff_daemon_CP_12469_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal RPIPE_w_out_buf_13993_inst_req_1 : boolean;
  signal RPIPE_w_out_buf_13993_inst_ack_1 : boolean;
  signal do_while_stmt_13990_branch_req_0 : boolean;
  signal RPIPE_w_out_buf_13993_inst_req_0 : boolean;
  signal RPIPE_w_out_buf_13993_inst_ack_0 : boolean;
  signal do_while_stmt_13990_branch_ack_1 : boolean;
  signal do_while_stmt_13990_branch_ack_0 : boolean;
  signal WPIPE_out_data_14006_inst_req_1 : boolean;
  signal WPIPE_out_data_14006_inst_ack_1 : boolean;
  signal WPIPE_out_data_14006_inst_req_0 : boolean;
  signal WPIPE_out_data_14006_inst_ack_0 : boolean;
  signal WPIPE_out_data_14003_inst_req_1 : boolean;
  signal WPIPE_out_data_14003_inst_ack_1 : boolean;
  signal WPIPE_out_data_14003_inst_req_0 : boolean;
  signal WPIPE_out_data_14003_inst_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "w_out_buff_daemon_input_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      bypass_flag => true,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  w_out_buff_daemon_CP_12469_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "w_out_buff_daemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= w_out_buff_daemon_CP_12469_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= w_out_buff_daemon_CP_12469_start & tag_ilock_write_ack_symbol;
    gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= w_out_buff_daemon_CP_12469_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  w_out_buff_daemon_CP_12469: Block -- control-path 
    signal w_out_buff_daemon_CP_12469_elements: BooleanArray(31 downto 0);
    -- 
  begin -- 
    w_out_buff_daemon_CP_12469_elements(0) <= w_out_buff_daemon_CP_12469_start;
    w_out_buff_daemon_CP_12469_symbol <= w_out_buff_daemon_CP_12469_elements(31);
    -- CP-element group 0:  transition  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (2) 
      -- CP-element group 0: 	 branch_block_stmt_13989/$entry
      -- CP-element group 0: 	 $entry
      -- 
    -- CP-element group 1:  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	3 
    -- CP-element group 1:  members (2) 
      -- CP-element group 1: 	 branch_block_stmt_13989/branch_block_stmt_13989__entry__
      -- CP-element group 1: 	 branch_block_stmt_13989/do_while_stmt_13990__entry__
      -- 
    w_out_buff_daemon_CP_12469_elements(1) <= w_out_buff_daemon_CP_12469_elements(0);
    -- CP-element group 2:  place  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	30 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	31 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_13989/branch_block_stmt_13989__exit__
      -- CP-element group 2: 	 branch_block_stmt_13989/do_while_stmt_13990__exit__
      -- 
    w_out_buff_daemon_CP_12469_elements(2) <= w_out_buff_daemon_CP_12469_elements(30);
    -- CP-element group 3:  transition  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	1 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_13989/do_while_stmt_13990/$entry
      -- 
    w_out_buff_daemon_CP_12469_elements(3) <= w_out_buff_daemon_CP_12469_elements(1);
    -- CP-element group 4:  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	10 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_13989/do_while_stmt_13990/do_while_stmt_13990__entry__
      -- 
    w_out_buff_daemon_CP_12469_elements(4) <= w_out_buff_daemon_CP_12469_elements(3);
    -- CP-element group 5:  merge  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	30 
    -- CP-element group 5:  members (1) 
      -- CP-element group 5: 	 branch_block_stmt_13989/do_while_stmt_13990/do_while_stmt_13990__exit__
      -- 
    -- Element group w_out_buff_daemon_CP_12469_elements(5) is bound as output of CP function.
    -- CP-element group 6:  merge  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	9 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_13989/do_while_stmt_13990/loop_back
      -- 
    -- Element group w_out_buff_daemon_CP_12469_elements(6) is bound as output of CP function.
    -- CP-element group 7:  branch  place  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	11 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	26 
    -- CP-element group 7: 	28 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_13989/do_while_stmt_13990/condition_done
      -- 
    w_out_buff_daemon_CP_12469_elements(7) <= w_out_buff_daemon_CP_12469_elements(11);
    -- CP-element group 8:  branch  place  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	25 
    -- CP-element group 8: successors 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_13989/do_while_stmt_13990/loop_body_done
      -- 
    w_out_buff_daemon_CP_12469_elements(8) <= w_out_buff_daemon_CP_12469_elements(25);
    -- CP-element group 9:  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	6 
    -- CP-element group 9: successors 
    -- CP-element group 9:  members (1) 
      -- CP-element group 9: 	 branch_block_stmt_13989/do_while_stmt_13990/do_while_stmt_13990_loop_body/back_edge_to_loop_body
      -- 
    w_out_buff_daemon_CP_12469_elements(9) <= w_out_buff_daemon_CP_12469_elements(6);
    -- CP-element group 10:  transition  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	4 
    -- CP-element group 10: successors 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_13989/do_while_stmt_13990/do_while_stmt_13990_loop_body/first_time_through_loop_body
      -- 
    w_out_buff_daemon_CP_12469_elements(10) <= w_out_buff_daemon_CP_12469_elements(4);
    -- CP-element group 11:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11: 	7 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 branch_block_stmt_13989/do_while_stmt_13990/do_while_stmt_13990_loop_body/loop_body_start
      -- CP-element group 11: 	 branch_block_stmt_13989/do_while_stmt_13990/do_while_stmt_13990_loop_body/condition_evaluated
      -- CP-element group 11: 	 branch_block_stmt_13989/do_while_stmt_13990/do_while_stmt_13990_loop_body/$entry
      -- 
    condition_evaluated_12493_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_12493_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => w_out_buff_daemon_CP_12469_elements(11), ack => do_while_stmt_13990_branch_req_0); -- 
    -- Element group w_out_buff_daemon_CP_12469_elements(11) is bound as output of CP function.
    -- CP-element group 12:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: marked-predecessors 
    -- CP-element group 12: 	14 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	14 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_13989/do_while_stmt_13990/do_while_stmt_13990_loop_body/RPIPE_w_out_buf_13993_sample_start_
      -- CP-element group 12: 	 branch_block_stmt_13989/do_while_stmt_13990/do_while_stmt_13990_loop_body/RPIPE_w_out_buf_13993_Sample/$entry
      -- CP-element group 12: 	 branch_block_stmt_13989/do_while_stmt_13990/do_while_stmt_13990_loop_body/RPIPE_w_out_buf_13993_Sample/rr
      -- 
    rr_12502_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_12502_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => w_out_buff_daemon_CP_12469_elements(12), ack => RPIPE_w_out_buf_13993_inst_req_0); -- 
    w_out_buff_daemon_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 37) := "w_out_buff_daemon_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= w_out_buff_daemon_CP_12469_elements(11) & w_out_buff_daemon_CP_12469_elements(14);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => w_out_buff_daemon_CP_12469_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	14 
    -- CP-element group 13: marked-predecessors 
    -- CP-element group 13: 	22 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	15 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 branch_block_stmt_13989/do_while_stmt_13990/do_while_stmt_13990_loop_body/RPIPE_w_out_buf_13993_Update/$entry
      -- CP-element group 13: 	 branch_block_stmt_13989/do_while_stmt_13990/do_while_stmt_13990_loop_body/RPIPE_w_out_buf_13993_Update/cr
      -- CP-element group 13: 	 branch_block_stmt_13989/do_while_stmt_13990/do_while_stmt_13990_loop_body/RPIPE_w_out_buf_13993_update_start_
      -- 
    cr_12507_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_12507_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => w_out_buff_daemon_CP_12469_elements(13), ack => RPIPE_w_out_buf_13993_inst_req_1); -- 
    w_out_buff_daemon_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "w_out_buff_daemon_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= w_out_buff_daemon_CP_12469_elements(14) & w_out_buff_daemon_CP_12469_elements(22);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => w_out_buff_daemon_CP_12469_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	12 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	12 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_13989/do_while_stmt_13990/do_while_stmt_13990_loop_body/RPIPE_w_out_buf_13993_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_13989/do_while_stmt_13990/do_while_stmt_13990_loop_body/RPIPE_w_out_buf_13993_Sample/$exit
      -- CP-element group 14: 	 branch_block_stmt_13989/do_while_stmt_13990/do_while_stmt_13990_loop_body/RPIPE_w_out_buf_13993_Sample/ra
      -- 
    ra_12503_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_w_out_buf_13993_inst_ack_0, ack => w_out_buff_daemon_CP_12469_elements(14)); -- 
    -- CP-element group 15:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	13 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15: 	20 
    -- CP-element group 15:  members (43) 
      -- CP-element group 15: 	 branch_block_stmt_13989/do_while_stmt_13990/do_while_stmt_13990_loop_body/RPIPE_w_out_buf_13993_Update/$exit
      -- CP-element group 15: 	 branch_block_stmt_13989/do_while_stmt_13990/do_while_stmt_13990_loop_body/RPIPE_w_out_buf_13993_Update/ca
      -- CP-element group 15: 	 branch_block_stmt_13989/do_while_stmt_13990/do_while_stmt_13990_loop_body/slice_13997_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_13989/do_while_stmt_13990/do_while_stmt_13990_loop_body/slice_13997_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_13989/do_while_stmt_13990/do_while_stmt_13990_loop_body/slice_13997_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_13989/do_while_stmt_13990/do_while_stmt_13990_loop_body/slice_13997_Sample/ra
      -- CP-element group 15: 	 branch_block_stmt_13989/do_while_stmt_13990/do_while_stmt_13990_loop_body/R_Z_13996_update_start_
      -- CP-element group 15: 	 branch_block_stmt_13989/do_while_stmt_13990/do_while_stmt_13990_loop_body/R_Z_13996_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_13989/do_while_stmt_13990/do_while_stmt_13990_loop_body/slice_13997_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_13989/do_while_stmt_13990/do_while_stmt_13990_loop_body/slice_13997_update_start_
      -- CP-element group 15: 	 branch_block_stmt_13989/do_while_stmt_13990/do_while_stmt_13990_loop_body/slice_13997_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_13989/do_while_stmt_13990/do_while_stmt_13990_loop_body/R_Z_13996_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_13989/do_while_stmt_13990/do_while_stmt_13990_loop_body/R_Z_13996_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_13989/do_while_stmt_13990/do_while_stmt_13990_loop_body/slice_13997_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_13989/do_while_stmt_13990/do_while_stmt_13990_loop_body/slice_13997_Update/$exit
      -- CP-element group 15: 	 branch_block_stmt_13989/do_while_stmt_13990/do_while_stmt_13990_loop_body/slice_13997_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_13989/do_while_stmt_13990/do_while_stmt_13990_loop_body/slice_13997_Update/ca
      -- CP-element group 15: 	 branch_block_stmt_13989/do_while_stmt_13990/do_while_stmt_13990_loop_body/RPIPE_w_out_buf_13993_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_13989/do_while_stmt_13990/do_while_stmt_13990_loop_body/slice_13997_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_13989/do_while_stmt_13990/do_while_stmt_13990_loop_body/R_Yb_14007_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_13989/do_while_stmt_13990/do_while_stmt_13990_loop_body/R_Yb_14007_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_13989/do_while_stmt_13990/do_while_stmt_13990_loop_body/R_Yb_14007_update_start_
      -- CP-element group 15: 	 branch_block_stmt_13989/do_while_stmt_13990/do_while_stmt_13990_loop_body/R_Yb_14007_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_13989/do_while_stmt_13990/do_while_stmt_13990_loop_body/R_Ya_14004_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_13989/do_while_stmt_13990/do_while_stmt_13990_loop_body/R_Ya_14004_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_13989/do_while_stmt_13990/do_while_stmt_13990_loop_body/R_Ya_14004_update_start_
      -- CP-element group 15: 	 branch_block_stmt_13989/do_while_stmt_13990/do_while_stmt_13990_loop_body/R_Ya_14004_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_13989/do_while_stmt_13990/do_while_stmt_13990_loop_body/slice_14001_Update/$exit
      -- CP-element group 15: 	 branch_block_stmt_13989/do_while_stmt_13990/do_while_stmt_13990_loop_body/slice_14001_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_13989/do_while_stmt_13990/do_while_stmt_13990_loop_body/slice_14001_Update/ca
      -- CP-element group 15: 	 branch_block_stmt_13989/do_while_stmt_13990/do_while_stmt_13990_loop_body/slice_14001_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_13989/do_while_stmt_13990/do_while_stmt_13990_loop_body/slice_14001_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_13989/do_while_stmt_13990/do_while_stmt_13990_loop_body/slice_14001_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_13989/do_while_stmt_13990/do_while_stmt_13990_loop_body/slice_14001_Sample/ra
      -- CP-element group 15: 	 branch_block_stmt_13989/do_while_stmt_13990/do_while_stmt_13990_loop_body/slice_14001_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_13989/do_while_stmt_13990/do_while_stmt_13990_loop_body/R_Z_14000_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_13989/do_while_stmt_13990/do_while_stmt_13990_loop_body/R_Z_14000_update_start_
      -- CP-element group 15: 	 branch_block_stmt_13989/do_while_stmt_13990/do_while_stmt_13990_loop_body/R_Z_14000_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_13989/do_while_stmt_13990/do_while_stmt_13990_loop_body/slice_14001_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_13989/do_while_stmt_13990/do_while_stmt_13990_loop_body/slice_14001_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_13989/do_while_stmt_13990/do_while_stmt_13990_loop_body/slice_14001_update_start_
      -- CP-element group 15: 	 branch_block_stmt_13989/do_while_stmt_13990/do_while_stmt_13990_loop_body/slice_14001_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_13989/do_while_stmt_13990/do_while_stmt_13990_loop_body/R_Z_14000_sample_start_
      -- 
    ca_12508_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_w_out_buf_13993_inst_ack_1, ack => w_out_buff_daemon_CP_12469_elements(15)); -- 
    -- CP-element group 16:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	22 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	18 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_13989/do_while_stmt_13990/do_while_stmt_13990_loop_body/WPIPE_out_data_14003_Sample/req
      -- CP-element group 16: 	 branch_block_stmt_13989/do_while_stmt_13990/do_while_stmt_13990_loop_body/WPIPE_out_data_14003_sample_start_
      -- CP-element group 16: 	 branch_block_stmt_13989/do_while_stmt_13990/do_while_stmt_13990_loop_body/WPIPE_out_data_14003_Sample/$entry
      -- 
    req_12556_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_12556_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => w_out_buff_daemon_CP_12469_elements(16), ack => WPIPE_out_data_14003_inst_req_0); -- 
    w_out_buff_daemon_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 37) := "w_out_buff_daemon_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= w_out_buff_daemon_CP_12469_elements(15) & w_out_buff_daemon_CP_12469_elements(22);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => w_out_buff_daemon_CP_12469_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	18 
    -- CP-element group 17: marked-predecessors 
    -- CP-element group 17: 	19 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	19 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 branch_block_stmt_13989/do_while_stmt_13990/do_while_stmt_13990_loop_body/WPIPE_out_data_14003_Update/req
      -- CP-element group 17: 	 branch_block_stmt_13989/do_while_stmt_13990/do_while_stmt_13990_loop_body/WPIPE_out_data_14003_Update/$entry
      -- CP-element group 17: 	 branch_block_stmt_13989/do_while_stmt_13990/do_while_stmt_13990_loop_body/WPIPE_out_data_14003_update_start_
      -- 
    req_12561_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_12561_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => w_out_buff_daemon_CP_12469_elements(17), ack => WPIPE_out_data_14003_inst_req_1); -- 
    w_out_buff_daemon_cp_element_group_17: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "w_out_buff_daemon_cp_element_group_17"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= w_out_buff_daemon_CP_12469_elements(18) & w_out_buff_daemon_CP_12469_elements(19);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => w_out_buff_daemon_CP_12469_elements(17), clk => clk, reset => reset); --
    end block;
    -- CP-element group 18:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	16 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: 	24 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 branch_block_stmt_13989/do_while_stmt_13990/do_while_stmt_13990_loop_body/WPIPE_out_data_14003_Sample/$exit
      -- CP-element group 18: 	 branch_block_stmt_13989/do_while_stmt_13990/do_while_stmt_13990_loop_body/WPIPE_out_data_14003_Sample/ack
      -- CP-element group 18: 	 branch_block_stmt_13989/do_while_stmt_13990/do_while_stmt_13990_loop_body/WPIPE_out_data_14003_sample_completed_
      -- 
    ack_12557_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_out_data_14003_inst_ack_0, ack => w_out_buff_daemon_CP_12469_elements(18)); -- 
    -- CP-element group 19:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	17 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	25 
    -- CP-element group 19: marked-successors 
    -- CP-element group 19: 	17 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_13989/do_while_stmt_13990/do_while_stmt_13990_loop_body/WPIPE_out_data_14003_Update/ack
      -- CP-element group 19: 	 branch_block_stmt_13989/do_while_stmt_13990/do_while_stmt_13990_loop_body/WPIPE_out_data_14003_Update/$exit
      -- CP-element group 19: 	 branch_block_stmt_13989/do_while_stmt_13990/do_while_stmt_13990_loop_body/WPIPE_out_data_14003_update_completed_
      -- 
    ack_12562_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_out_data_14003_inst_ack_1, ack => w_out_buff_daemon_CP_12469_elements(19)); -- 
    -- CP-element group 20:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	15 
    -- CP-element group 20: 	24 
    -- CP-element group 20: marked-predecessors 
    -- CP-element group 20: 	22 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	22 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_13989/do_while_stmt_13990/do_while_stmt_13990_loop_body/WPIPE_out_data_14006_Sample/$entry
      -- CP-element group 20: 	 branch_block_stmt_13989/do_while_stmt_13990/do_while_stmt_13990_loop_body/WPIPE_out_data_14006_Sample/req
      -- CP-element group 20: 	 branch_block_stmt_13989/do_while_stmt_13990/do_while_stmt_13990_loop_body/WPIPE_out_data_14006_sample_start_
      -- 
    req_12574_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_12574_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => w_out_buff_daemon_CP_12469_elements(20), ack => WPIPE_out_data_14006_inst_req_0); -- 
    w_out_buff_daemon_cp_element_group_20: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 3,1 => 3,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 37) := "w_out_buff_daemon_cp_element_group_20"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= w_out_buff_daemon_CP_12469_elements(15) & w_out_buff_daemon_CP_12469_elements(24) & w_out_buff_daemon_CP_12469_elements(22);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => w_out_buff_daemon_CP_12469_elements(20), clk => clk, reset => reset); --
    end block;
    -- CP-element group 21:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	22 
    -- CP-element group 21: marked-predecessors 
    -- CP-element group 21: 	23 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	23 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_13989/do_while_stmt_13990/do_while_stmt_13990_loop_body/WPIPE_out_data_14006_Update/req
      -- CP-element group 21: 	 branch_block_stmt_13989/do_while_stmt_13990/do_while_stmt_13990_loop_body/WPIPE_out_data_14006_Update/$entry
      -- CP-element group 21: 	 branch_block_stmt_13989/do_while_stmt_13990/do_while_stmt_13990_loop_body/WPIPE_out_data_14006_update_start_
      -- 
    req_12579_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_12579_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => w_out_buff_daemon_CP_12469_elements(21), ack => WPIPE_out_data_14006_inst_req_1); -- 
    w_out_buff_daemon_cp_element_group_21: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "w_out_buff_daemon_cp_element_group_21"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= w_out_buff_daemon_CP_12469_elements(22) & w_out_buff_daemon_CP_12469_elements(23);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => w_out_buff_daemon_CP_12469_elements(21), clk => clk, reset => reset); --
    end block;
    -- CP-element group 22:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	20 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: marked-successors 
    -- CP-element group 22: 	16 
    -- CP-element group 22: 	20 
    -- CP-element group 22: 	13 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_13989/do_while_stmt_13990/do_while_stmt_13990_loop_body/WPIPE_out_data_14006_Sample/$exit
      -- CP-element group 22: 	 branch_block_stmt_13989/do_while_stmt_13990/do_while_stmt_13990_loop_body/WPIPE_out_data_14006_Sample/ack
      -- CP-element group 22: 	 branch_block_stmt_13989/do_while_stmt_13990/do_while_stmt_13990_loop_body/WPIPE_out_data_14006_sample_completed_
      -- 
    ack_12575_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_out_data_14006_inst_ack_0, ack => w_out_buff_daemon_CP_12469_elements(22)); -- 
    -- CP-element group 23:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	21 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	25 
    -- CP-element group 23: marked-successors 
    -- CP-element group 23: 	21 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_13989/do_while_stmt_13990/do_while_stmt_13990_loop_body/WPIPE_out_data_14006_Update/$exit
      -- CP-element group 23: 	 branch_block_stmt_13989/do_while_stmt_13990/do_while_stmt_13990_loop_body/WPIPE_out_data_14006_Update/ack
      -- CP-element group 23: 	 branch_block_stmt_13989/do_while_stmt_13990/do_while_stmt_13990_loop_body/WPIPE_out_data_14006_update_completed_
      -- 
    ack_12580_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_out_data_14006_inst_ack_1, ack => w_out_buff_daemon_CP_12469_elements(23)); -- 
    -- CP-element group 24:  transition  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	18 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	20 
    -- CP-element group 24:  members (1) 
      -- CP-element group 24: 	 branch_block_stmt_13989/do_while_stmt_13990/do_while_stmt_13990_loop_body/delay_transition_14003_14006
      -- 
    -- Element group w_out_buff_daemon_CP_12469_elements(24) is a control-delay.
    cp_element_24_delay: control_delay_element  generic map(name => " 24_delay", delay_value => 1)  port map(req => w_out_buff_daemon_CP_12469_elements(18), ack => w_out_buff_daemon_CP_12469_elements(24), clk => clk, reset =>reset);
    -- CP-element group 25:  join  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	23 
    -- CP-element group 25: 	19 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	8 
    -- CP-element group 25:  members (1) 
      -- CP-element group 25: 	 branch_block_stmt_13989/do_while_stmt_13990/do_while_stmt_13990_loop_body/$exit
      -- 
    w_out_buff_daemon_cp_element_group_25: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 3);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "w_out_buff_daemon_cp_element_group_25"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= w_out_buff_daemon_CP_12469_elements(23) & w_out_buff_daemon_CP_12469_elements(19);
      gj : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => w_out_buff_daemon_CP_12469_elements(25), clk => clk, reset => reset); --
    end block;
    -- CP-element group 26:  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	7 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	27 
    -- CP-element group 26:  members (1) 
      -- CP-element group 26: 	 branch_block_stmt_13989/do_while_stmt_13990/loop_exit/$entry
      -- 
    w_out_buff_daemon_CP_12469_elements(26) <= w_out_buff_daemon_CP_12469_elements(7);
    -- CP-element group 27:  transition  input  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	26 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (2) 
      -- CP-element group 27: 	 branch_block_stmt_13989/do_while_stmt_13990/loop_exit/$exit
      -- CP-element group 27: 	 branch_block_stmt_13989/do_while_stmt_13990/loop_exit/ack
      -- 
    ack_12585_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_13990_branch_ack_0, ack => w_out_buff_daemon_CP_12469_elements(27)); -- 
    -- CP-element group 28:  transition  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	7 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28:  members (1) 
      -- CP-element group 28: 	 branch_block_stmt_13989/do_while_stmt_13990/loop_taken/$entry
      -- 
    w_out_buff_daemon_CP_12469_elements(28) <= w_out_buff_daemon_CP_12469_elements(7);
    -- CP-element group 29:  transition  input  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	28 
    -- CP-element group 29: successors 
    -- CP-element group 29:  members (2) 
      -- CP-element group 29: 	 branch_block_stmt_13989/do_while_stmt_13990/loop_taken/ack
      -- CP-element group 29: 	 branch_block_stmt_13989/do_while_stmt_13990/loop_taken/$exit
      -- 
    ack_12589_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_13990_branch_ack_1, ack => w_out_buff_daemon_CP_12469_elements(29)); -- 
    -- CP-element group 30:  transition  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	5 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	2 
    -- CP-element group 30:  members (1) 
      -- CP-element group 30: 	 branch_block_stmt_13989/do_while_stmt_13990/$exit
      -- 
    w_out_buff_daemon_CP_12469_elements(30) <= w_out_buff_daemon_CP_12469_elements(5);
    -- CP-element group 31:  transition  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	2 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (2) 
      -- CP-element group 31: 	 branch_block_stmt_13989/$exit
      -- CP-element group 31: 	 $exit
      -- 
    w_out_buff_daemon_CP_12469_elements(31) <= w_out_buff_daemon_CP_12469_elements(2);
    do_while_stmt_13990_terminator_12590: loop_terminator -- 
      generic map (name => " do_while_stmt_13990_terminator_12590", max_iterations_in_flight =>3) 
      port map(loop_body_exit => w_out_buff_daemon_CP_12469_elements(8),loop_continue => w_out_buff_daemon_CP_12469_elements(29),loop_terminate => w_out_buff_daemon_CP_12469_elements(27),loop_back => w_out_buff_daemon_CP_12469_elements(6),loop_exit => w_out_buff_daemon_CP_12469_elements(5),clk => clk, reset => reset); -- 
    entry_tmerge_12494_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= w_out_buff_daemon_CP_12469_elements(9);
        preds(1)  <= w_out_buff_daemon_CP_12469_elements(10);
        entry_tmerge_12494 : transition_merge -- 
          generic map(name => " entry_tmerge_12494")
          port map (preds => preds, symbol_out => w_out_buff_daemon_CP_12469_elements(11));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal Ya_13998 : std_logic_vector(63 downto 0);
    signal Yb_14002 : std_logic_vector(63 downto 0);
    signal Z_13994 : std_logic_vector(127 downto 0);
    signal konst_14010_wire_constant : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    konst_14010_wire_constant <= "1";
    -- flow-through slice operator slice_13997_inst
    Ya_13998 <= Z_13994(127 downto 64);
    -- flow-through slice operator slice_14001_inst
    Yb_14002 <= Z_13994(63 downto 0);
    do_while_stmt_13990_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= konst_14010_wire_constant;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_13990_branch", condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_13990_branch_req_0,
          ack0 => do_while_stmt_13990_branch_ack_0,
          ack1 => do_while_stmt_13990_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- shared inport operator group (0) : RPIPE_w_out_buf_13993_inst 
    InportGroup0: Block -- 
      signal data_out: std_logic_vector(127 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_w_out_buf_13993_inst_req_0;
      RPIPE_w_out_buf_13993_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_w_out_buf_13993_inst_req_1;
      RPIPE_w_out_buf_13993_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      gI: SplitGuardInterface generic map(name => "gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Z_13994 <= data_out(127 downto 0);
      w_out_buf_read_0: InputPortRevised -- 
        generic map ( name => "w_out_buf_read_0", data_width => 128,  num_reqs => 1,  output_buffering => outBUFs,   no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => w_out_buf_pipe_read_req(0),
          oack => w_out_buf_pipe_read_ack(0),
          odata => w_out_buf_pipe_read_data(127 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_out_data_14006_inst WPIPE_out_data_14003_inst 
    OutportGroup0: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal sample_req, sample_ack : BooleanArray( 1 downto 0);
      signal update_req, update_ack : BooleanArray( 1 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 1 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      sample_req_unguarded(1) <= WPIPE_out_data_14006_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_out_data_14003_inst_req_0;
      WPIPE_out_data_14006_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_out_data_14003_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(1) <= WPIPE_out_data_14006_inst_req_1;
      update_req_unguarded(0) <= WPIPE_out_data_14003_inst_req_1;
      WPIPE_out_data_14006_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_out_data_14003_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      gI: SplitGuardInterface generic map(name => "gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      data_in <= Yb_14002 & Ya_13998;
      out_data_write_0: OutputPortRevised -- 
        generic map ( name => "out_data", data_width => 64, num_reqs => 2, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => out_data_pipe_write_req(0),
          oack => out_data_pipe_write_ack(0),
          odata => out_data_pipe_write_data(63 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end w_out_buff_daemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library work;
use work.ahir_system_global_package.all;
entity ahir_system is  -- system 
  port (-- 
    clk : in std_logic;
    reset : in std_logic;
    in_data_pipe_write_data: in std_logic_vector(63 downto 0);
    in_data_pipe_write_req : in std_logic_vector(0 downto 0);
    in_data_pipe_write_ack : out std_logic_vector(0 downto 0);
    out_data_pipe_read_data: out std_logic_vector(63 downto 0);
    out_data_pipe_read_req : in std_logic_vector(0 downto 0);
    out_data_pipe_read_ack : out std_logic_vector(0 downto 0)); -- 
  -- 
end entity; 
architecture ahir_system_arch  of ahir_system is -- system-architecture 
  -- declarations related to module In_wrap_daemon
  component In_wrap_daemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      w_in_buf_pipe_read_req : out  std_logic_vector(0 downto 0);
      w_in_buf_pipe_read_ack : in   std_logic_vector(0 downto 0);
      w_in_buf_pipe_read_data : in   std_logic_vector(127 downto 0);
      cmd_in_pipe_write_req : out  std_logic_vector(0 downto 0);
      cmd_in_pipe_write_ack : in   std_logic_vector(0 downto 0);
      cmd_in_pipe_write_data : out  std_logic_vector(63 downto 0);
      d_in_buf_pipe_write_req : out  std_logic_vector(0 downto 0);
      d_in_buf_pipe_write_ack : in   std_logic_vector(0 downto 0);
      d_in_buf_pipe_write_data : out  std_logic_vector(127 downto 0);
      e_in_buf_pipe_write_req : out  std_logic_vector(0 downto 0);
      e_in_buf_pipe_write_ack : in   std_logic_vector(0 downto 0);
      e_in_buf_pipe_write_data : out  std_logic_vector(127 downto 0);
      out_wrap_cmd_pipe_write_req : out  std_logic_vector(0 downto 0);
      out_wrap_cmd_pipe_write_ack : in   std_logic_vector(0 downto 0);
      out_wrap_cmd_pipe_write_data : out  std_logic_vector(63 downto 0);
      out_wrap_data_pipe_write_req : out  std_logic_vector(0 downto 0);
      out_wrap_data_pipe_write_ack : in   std_logic_vector(0 downto 0);
      out_wrap_data_pipe_write_data : out  std_logic_vector(127 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module In_wrap_daemon
  signal In_wrap_daemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal In_wrap_daemon_tag_out   : std_logic_vector(1 downto 0);
  signal In_wrap_daemon_start_req : std_logic;
  signal In_wrap_daemon_start_ack : std_logic;
  signal In_wrap_daemon_fin_req   : std_logic;
  signal In_wrap_daemon_fin_ack : std_logic;
  -- declarations related to module Inv_Sbox_1
  -- declarations related to module Inv_Sbox_2
  -- declarations related to module Inv_Sbox_3
  -- declarations related to module Inv_Sbox_4
  -- declarations related to module MUL2
  -- declarations related to module Out_wrap_daemon
  component Out_wrap_daemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      e_out_buf_pipe_read_req : out  std_logic_vector(0 downto 0);
      e_out_buf_pipe_read_ack : in   std_logic_vector(0 downto 0);
      e_out_buf_pipe_read_data : in   std_logic_vector(127 downto 0);
      d_out_buf_pipe_read_req : out  std_logic_vector(0 downto 0);
      d_out_buf_pipe_read_ack : in   std_logic_vector(0 downto 0);
      d_out_buf_pipe_read_data : in   std_logic_vector(127 downto 0);
      out_wrap_cmd_pipe_read_req : out  std_logic_vector(0 downto 0);
      out_wrap_cmd_pipe_read_ack : in   std_logic_vector(0 downto 0);
      out_wrap_cmd_pipe_read_data : in   std_logic_vector(63 downto 0);
      out_wrap_data_pipe_read_req : out  std_logic_vector(0 downto 0);
      out_wrap_data_pipe_read_ack : in   std_logic_vector(0 downto 0);
      out_wrap_data_pipe_read_data : in   std_logic_vector(127 downto 0);
      status_out_pipe_read_req : out  std_logic_vector(0 downto 0);
      status_out_pipe_read_ack : in   std_logic_vector(0 downto 0);
      status_out_pipe_read_data : in   std_logic_vector(63 downto 0);
      w_out_buf_pipe_write_req : out  std_logic_vector(0 downto 0);
      w_out_buf_pipe_write_ack : in   std_logic_vector(0 downto 0);
      w_out_buf_pipe_write_data : out  std_logic_vector(127 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module Out_wrap_daemon
  signal Out_wrap_daemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal Out_wrap_daemon_tag_out   : std_logic_vector(1 downto 0);
  signal Out_wrap_daemon_start_req : std_logic;
  signal Out_wrap_daemon_start_ack : std_logic;
  signal Out_wrap_daemon_fin_req   : std_logic;
  signal Out_wrap_daemon_fin_ack : std_logic;
  -- declarations related to module c_block_daemon
  component c_block_daemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      cmd_in_pipe_read_req : out  std_logic_vector(0 downto 0);
      cmd_in_pipe_read_ack : in   std_logic_vector(0 downto 0);
      cmd_in_pipe_read_data : in   std_logic_vector(63 downto 0);
      d_block_done_pipe_read_req : out  std_logic_vector(0 downto 0);
      d_block_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
      d_block_done_pipe_read_data : in   std_logic_vector(0 downto 0);
      e_block_done_pipe_read_req : out  std_logic_vector(0 downto 0);
      e_block_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
      e_block_done_pipe_read_data : in   std_logic_vector(0 downto 0);
      d_cmd_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      d_cmd_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      d_cmd_pipe_pipe_write_data : out  std_logic_vector(143 downto 0);
      e_cmd_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      e_cmd_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      e_cmd_pipe_pipe_write_data : out  std_logic_vector(143 downto 0);
      status_out_pipe_write_req : out  std_logic_vector(0 downto 0);
      status_out_pipe_write_ack : in   std_logic_vector(0 downto 0);
      status_out_pipe_write_data : out  std_logic_vector(63 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module c_block_daemon
  signal c_block_daemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal c_block_daemon_tag_out   : std_logic_vector(1 downto 0);
  signal c_block_daemon_start_req : std_logic;
  signal c_block_daemon_start_ack : std_logic;
  signal c_block_daemon_fin_req   : std_logic;
  signal c_block_daemon_fin_ack : std_logic;
  -- declarations related to module d_block_daemon
  component d_block_daemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      d_cmd_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      d_cmd_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      d_cmd_pipe_pipe_read_data : in   std_logic_vector(143 downto 0);
      d_in_buf_pipe_read_req : out  std_logic_vector(0 downto 0);
      d_in_buf_pipe_read_ack : in   std_logic_vector(0 downto 0);
      d_in_buf_pipe_read_data : in   std_logic_vector(127 downto 0);
      d_block_done_pipe_write_req : out  std_logic_vector(0 downto 0);
      d_block_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
      d_block_done_pipe_write_data : out  std_logic_vector(0 downto 0);
      d_out_buf_pipe_write_req : out  std_logic_vector(0 downto 0);
      d_out_buf_pipe_write_ack : in   std_logic_vector(0 downto 0);
      d_out_buf_pipe_write_data : out  std_logic_vector(127 downto 0);
      key_expand_single_call_reqs : out  std_logic_vector(0 downto 0);
      key_expand_single_call_acks : in   std_logic_vector(0 downto 0);
      key_expand_single_call_data : out  std_logic_vector(135 downto 0);
      key_expand_single_call_tag  :  out  std_logic_vector(3 downto 0);
      key_expand_single_return_reqs : out  std_logic_vector(0 downto 0);
      key_expand_single_return_acks : in   std_logic_vector(0 downto 0);
      key_expand_single_return_data : in   std_logic_vector(135 downto 0);
      key_expand_single_return_tag :  in   std_logic_vector(3 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module d_block_daemon
  signal d_block_daemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal d_block_daemon_tag_out   : std_logic_vector(1 downto 0);
  signal d_block_daemon_start_req : std_logic;
  signal d_block_daemon_start_ack : std_logic;
  signal d_block_daemon_fin_req   : std_logic;
  signal d_block_daemon_fin_ack : std_logic;
  -- declarations related to module dec_round
  -- declarations related to module e_block_daemon
  component e_block_daemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      e_in_buf_pipe_read_req : out  std_logic_vector(0 downto 0);
      e_in_buf_pipe_read_ack : in   std_logic_vector(0 downto 0);
      e_in_buf_pipe_read_data : in   std_logic_vector(127 downto 0);
      e_cmd_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      e_cmd_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      e_cmd_pipe_pipe_read_data : in   std_logic_vector(143 downto 0);
      e_out_buf_pipe_write_req : out  std_logic_vector(0 downto 0);
      e_out_buf_pipe_write_ack : in   std_logic_vector(0 downto 0);
      e_out_buf_pipe_write_data : out  std_logic_vector(127 downto 0);
      e_block_done_pipe_write_req : out  std_logic_vector(0 downto 0);
      e_block_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
      e_block_done_pipe_write_data : out  std_logic_vector(0 downto 0);
      key_expand_single_call_reqs : out  std_logic_vector(0 downto 0);
      key_expand_single_call_acks : in   std_logic_vector(0 downto 0);
      key_expand_single_call_data : out  std_logic_vector(135 downto 0);
      key_expand_single_call_tag  :  out  std_logic_vector(3 downto 0);
      key_expand_single_return_reqs : out  std_logic_vector(0 downto 0);
      key_expand_single_return_acks : in   std_logic_vector(0 downto 0);
      key_expand_single_return_data : in   std_logic_vector(135 downto 0);
      key_expand_single_return_tag :  in   std_logic_vector(3 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module e_block_daemon
  signal e_block_daemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal e_block_daemon_tag_out   : std_logic_vector(1 downto 0);
  signal e_block_daemon_start_req : std_logic;
  signal e_block_daemon_start_ack : std_logic;
  signal e_block_daemon_fin_req   : std_logic;
  signal e_block_daemon_fin_ack : std_logic;
  -- declarations related to module enc_round
  -- declarations related to module key_expand_single
  component key_expand_single is -- 
    generic (tag_length : integer); 
    port ( -- 
      K_in : in  std_logic_vector(127 downto 0);
      Round_C : in  std_logic_vector(7 downto 0);
      K_out : out  std_logic_vector(127 downto 0);
      nRound_C : out  std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module key_expand_single
  signal key_expand_single_K_in :  std_logic_vector(127 downto 0);
  signal key_expand_single_Round_C :  std_logic_vector(7 downto 0);
  signal key_expand_single_K_out :  std_logic_vector(127 downto 0);
  signal key_expand_single_nRound_C :  std_logic_vector(7 downto 0);
  signal key_expand_single_in_args    : std_logic_vector(135 downto 0);
  signal key_expand_single_out_args   : std_logic_vector(135 downto 0);
  signal key_expand_single_tag_in    : std_logic_vector(5 downto 0) := (others => '0');
  signal key_expand_single_tag_out   : std_logic_vector(5 downto 0);
  signal key_expand_single_start_req : std_logic;
  signal key_expand_single_start_ack : std_logic;
  signal key_expand_single_fin_req   : std_logic;
  signal key_expand_single_fin_ack : std_logic;
  -- caller side aggregated signals for module key_expand_single
  signal key_expand_single_call_reqs: std_logic_vector(1 downto 0);
  signal key_expand_single_call_acks: std_logic_vector(1 downto 0);
  signal key_expand_single_return_reqs: std_logic_vector(1 downto 0);
  signal key_expand_single_return_acks: std_logic_vector(1 downto 0);
  signal key_expand_single_call_data: std_logic_vector(271 downto 0);
  signal key_expand_single_call_tag: std_logic_vector(7 downto 0);
  signal key_expand_single_return_data: std_logic_vector(271 downto 0);
  signal key_expand_single_return_tag: std_logic_vector(7 downto 0);
  -- declarations related to module sbox_mux_impl
  -- declarations related to module w_in_buff_daemon
  component w_in_buff_daemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      in_data_pipe_read_req : out  std_logic_vector(0 downto 0);
      in_data_pipe_read_ack : in   std_logic_vector(0 downto 0);
      in_data_pipe_read_data : in   std_logic_vector(63 downto 0);
      w_in_buf_pipe_write_req : out  std_logic_vector(0 downto 0);
      w_in_buf_pipe_write_ack : in   std_logic_vector(0 downto 0);
      w_in_buf_pipe_write_data : out  std_logic_vector(127 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module w_in_buff_daemon
  signal w_in_buff_daemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal w_in_buff_daemon_tag_out   : std_logic_vector(1 downto 0);
  signal w_in_buff_daemon_start_req : std_logic;
  signal w_in_buff_daemon_start_ack : std_logic;
  signal w_in_buff_daemon_fin_req   : std_logic;
  signal w_in_buff_daemon_fin_ack : std_logic;
  -- declarations related to module w_out_buff_daemon
  component w_out_buff_daemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      w_out_buf_pipe_read_req : out  std_logic_vector(0 downto 0);
      w_out_buf_pipe_read_ack : in   std_logic_vector(0 downto 0);
      w_out_buf_pipe_read_data : in   std_logic_vector(127 downto 0);
      out_data_pipe_write_req : out  std_logic_vector(0 downto 0);
      out_data_pipe_write_ack : in   std_logic_vector(0 downto 0);
      out_data_pipe_write_data : out  std_logic_vector(63 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module w_out_buff_daemon
  signal w_out_buff_daemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal w_out_buff_daemon_tag_out   : std_logic_vector(1 downto 0);
  signal w_out_buff_daemon_start_req : std_logic;
  signal w_out_buff_daemon_start_ack : std_logic;
  signal w_out_buff_daemon_fin_req   : std_logic;
  signal w_out_buff_daemon_fin_ack : std_logic;
  -- aggregate signals for write to pipe cmd_in
  signal cmd_in_pipe_write_data: std_logic_vector(63 downto 0);
  signal cmd_in_pipe_write_req: std_logic_vector(0 downto 0);
  signal cmd_in_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe cmd_in
  signal cmd_in_pipe_read_data: std_logic_vector(63 downto 0);
  signal cmd_in_pipe_read_req: std_logic_vector(0 downto 0);
  signal cmd_in_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe d_block_done
  signal d_block_done_pipe_write_data: std_logic_vector(0 downto 0);
  signal d_block_done_pipe_write_req: std_logic_vector(0 downto 0);
  signal d_block_done_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe d_block_done
  signal d_block_done_pipe_read_data: std_logic_vector(0 downto 0);
  signal d_block_done_pipe_read_req: std_logic_vector(0 downto 0);
  signal d_block_done_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe d_cmd_pipe
  signal d_cmd_pipe_pipe_write_data: std_logic_vector(143 downto 0);
  signal d_cmd_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal d_cmd_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe d_cmd_pipe
  signal d_cmd_pipe_pipe_read_data: std_logic_vector(143 downto 0);
  signal d_cmd_pipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal d_cmd_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe d_in_buf
  signal d_in_buf_pipe_write_data: std_logic_vector(127 downto 0);
  signal d_in_buf_pipe_write_req: std_logic_vector(0 downto 0);
  signal d_in_buf_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe d_in_buf
  signal d_in_buf_pipe_read_data: std_logic_vector(127 downto 0);
  signal d_in_buf_pipe_read_req: std_logic_vector(0 downto 0);
  signal d_in_buf_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe d_out_buf
  signal d_out_buf_pipe_write_data: std_logic_vector(127 downto 0);
  signal d_out_buf_pipe_write_req: std_logic_vector(0 downto 0);
  signal d_out_buf_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe d_out_buf
  signal d_out_buf_pipe_read_data: std_logic_vector(127 downto 0);
  signal d_out_buf_pipe_read_req: std_logic_vector(0 downto 0);
  signal d_out_buf_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe e_block_done
  signal e_block_done_pipe_write_data: std_logic_vector(0 downto 0);
  signal e_block_done_pipe_write_req: std_logic_vector(0 downto 0);
  signal e_block_done_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe e_block_done
  signal e_block_done_pipe_read_data: std_logic_vector(0 downto 0);
  signal e_block_done_pipe_read_req: std_logic_vector(0 downto 0);
  signal e_block_done_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe e_cmd_pipe
  signal e_cmd_pipe_pipe_write_data: std_logic_vector(143 downto 0);
  signal e_cmd_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal e_cmd_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe e_cmd_pipe
  signal e_cmd_pipe_pipe_read_data: std_logic_vector(143 downto 0);
  signal e_cmd_pipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal e_cmd_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe e_in_buf
  signal e_in_buf_pipe_write_data: std_logic_vector(127 downto 0);
  signal e_in_buf_pipe_write_req: std_logic_vector(0 downto 0);
  signal e_in_buf_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe e_in_buf
  signal e_in_buf_pipe_read_data: std_logic_vector(127 downto 0);
  signal e_in_buf_pipe_read_req: std_logic_vector(0 downto 0);
  signal e_in_buf_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe e_out_buf
  signal e_out_buf_pipe_write_data: std_logic_vector(127 downto 0);
  signal e_out_buf_pipe_write_req: std_logic_vector(0 downto 0);
  signal e_out_buf_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe e_out_buf
  signal e_out_buf_pipe_read_data: std_logic_vector(127 downto 0);
  signal e_out_buf_pipe_read_req: std_logic_vector(0 downto 0);
  signal e_out_buf_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe in_data
  signal in_data_pipe_read_data: std_logic_vector(63 downto 0);
  signal in_data_pipe_read_req: std_logic_vector(0 downto 0);
  signal in_data_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe out_data
  signal out_data_pipe_write_data: std_logic_vector(63 downto 0);
  signal out_data_pipe_write_req: std_logic_vector(0 downto 0);
  signal out_data_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe out_wrap_cmd
  signal out_wrap_cmd_pipe_write_data: std_logic_vector(63 downto 0);
  signal out_wrap_cmd_pipe_write_req: std_logic_vector(0 downto 0);
  signal out_wrap_cmd_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe out_wrap_cmd
  signal out_wrap_cmd_pipe_read_data: std_logic_vector(63 downto 0);
  signal out_wrap_cmd_pipe_read_req: std_logic_vector(0 downto 0);
  signal out_wrap_cmd_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe out_wrap_data
  signal out_wrap_data_pipe_write_data: std_logic_vector(127 downto 0);
  signal out_wrap_data_pipe_write_req: std_logic_vector(0 downto 0);
  signal out_wrap_data_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe out_wrap_data
  signal out_wrap_data_pipe_read_data: std_logic_vector(127 downto 0);
  signal out_wrap_data_pipe_read_req: std_logic_vector(0 downto 0);
  signal out_wrap_data_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe status_out
  signal status_out_pipe_write_data: std_logic_vector(63 downto 0);
  signal status_out_pipe_write_req: std_logic_vector(0 downto 0);
  signal status_out_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe status_out
  signal status_out_pipe_read_data: std_logic_vector(63 downto 0);
  signal status_out_pipe_read_req: std_logic_vector(0 downto 0);
  signal status_out_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe w_in_buf
  signal w_in_buf_pipe_write_data: std_logic_vector(127 downto 0);
  signal w_in_buf_pipe_write_req: std_logic_vector(0 downto 0);
  signal w_in_buf_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe w_in_buf
  signal w_in_buf_pipe_read_data: std_logic_vector(127 downto 0);
  signal w_in_buf_pipe_read_req: std_logic_vector(0 downto 0);
  signal w_in_buf_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe w_out_buf
  signal w_out_buf_pipe_write_data: std_logic_vector(127 downto 0);
  signal w_out_buf_pipe_write_req: std_logic_vector(0 downto 0);
  signal w_out_buf_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe w_out_buf
  signal w_out_buf_pipe_read_data: std_logic_vector(127 downto 0);
  signal w_out_buf_pipe_read_req: std_logic_vector(0 downto 0);
  signal w_out_buf_pipe_read_ack: std_logic_vector(0 downto 0);
  -- 
begin -- 
  -- module In_wrap_daemon
  In_wrap_daemon_instance:In_wrap_daemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => In_wrap_daemon_start_req,
      start_ack => In_wrap_daemon_start_ack,
      fin_req => In_wrap_daemon_fin_req,
      fin_ack => In_wrap_daemon_fin_ack,
      clk => clk,
      reset => reset,
      w_in_buf_pipe_read_req => w_in_buf_pipe_read_req(0 downto 0),
      w_in_buf_pipe_read_ack => w_in_buf_pipe_read_ack(0 downto 0),
      w_in_buf_pipe_read_data => w_in_buf_pipe_read_data(127 downto 0),
      cmd_in_pipe_write_req => cmd_in_pipe_write_req(0 downto 0),
      cmd_in_pipe_write_ack => cmd_in_pipe_write_ack(0 downto 0),
      cmd_in_pipe_write_data => cmd_in_pipe_write_data(63 downto 0),
      d_in_buf_pipe_write_req => d_in_buf_pipe_write_req(0 downto 0),
      d_in_buf_pipe_write_ack => d_in_buf_pipe_write_ack(0 downto 0),
      d_in_buf_pipe_write_data => d_in_buf_pipe_write_data(127 downto 0),
      e_in_buf_pipe_write_req => e_in_buf_pipe_write_req(0 downto 0),
      e_in_buf_pipe_write_ack => e_in_buf_pipe_write_ack(0 downto 0),
      e_in_buf_pipe_write_data => e_in_buf_pipe_write_data(127 downto 0),
      out_wrap_cmd_pipe_write_req => out_wrap_cmd_pipe_write_req(0 downto 0),
      out_wrap_cmd_pipe_write_ack => out_wrap_cmd_pipe_write_ack(0 downto 0),
      out_wrap_cmd_pipe_write_data => out_wrap_cmd_pipe_write_data(63 downto 0),
      out_wrap_data_pipe_write_req => out_wrap_data_pipe_write_req(0 downto 0),
      out_wrap_data_pipe_write_ack => out_wrap_data_pipe_write_ack(0 downto 0),
      out_wrap_data_pipe_write_data => out_wrap_data_pipe_write_data(127 downto 0),
      tag_in => In_wrap_daemon_tag_in,
      tag_out => In_wrap_daemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  In_wrap_daemon_tag_in <= (others => '0');
  In_wrap_daemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => In_wrap_daemon_start_req, start_ack => In_wrap_daemon_start_ack,  fin_req => In_wrap_daemon_fin_req,  fin_ack => In_wrap_daemon_fin_ack);
  -- module Out_wrap_daemon
  Out_wrap_daemon_instance:Out_wrap_daemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => Out_wrap_daemon_start_req,
      start_ack => Out_wrap_daemon_start_ack,
      fin_req => Out_wrap_daemon_fin_req,
      fin_ack => Out_wrap_daemon_fin_ack,
      clk => clk,
      reset => reset,
      e_out_buf_pipe_read_req => e_out_buf_pipe_read_req(0 downto 0),
      e_out_buf_pipe_read_ack => e_out_buf_pipe_read_ack(0 downto 0),
      e_out_buf_pipe_read_data => e_out_buf_pipe_read_data(127 downto 0),
      d_out_buf_pipe_read_req => d_out_buf_pipe_read_req(0 downto 0),
      d_out_buf_pipe_read_ack => d_out_buf_pipe_read_ack(0 downto 0),
      d_out_buf_pipe_read_data => d_out_buf_pipe_read_data(127 downto 0),
      out_wrap_cmd_pipe_read_req => out_wrap_cmd_pipe_read_req(0 downto 0),
      out_wrap_cmd_pipe_read_ack => out_wrap_cmd_pipe_read_ack(0 downto 0),
      out_wrap_cmd_pipe_read_data => out_wrap_cmd_pipe_read_data(63 downto 0),
      out_wrap_data_pipe_read_req => out_wrap_data_pipe_read_req(0 downto 0),
      out_wrap_data_pipe_read_ack => out_wrap_data_pipe_read_ack(0 downto 0),
      out_wrap_data_pipe_read_data => out_wrap_data_pipe_read_data(127 downto 0),
      status_out_pipe_read_req => status_out_pipe_read_req(0 downto 0),
      status_out_pipe_read_ack => status_out_pipe_read_ack(0 downto 0),
      status_out_pipe_read_data => status_out_pipe_read_data(63 downto 0),
      w_out_buf_pipe_write_req => w_out_buf_pipe_write_req(0 downto 0),
      w_out_buf_pipe_write_ack => w_out_buf_pipe_write_ack(0 downto 0),
      w_out_buf_pipe_write_data => w_out_buf_pipe_write_data(127 downto 0),
      tag_in => Out_wrap_daemon_tag_in,
      tag_out => Out_wrap_daemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  Out_wrap_daemon_tag_in <= (others => '0');
  Out_wrap_daemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => Out_wrap_daemon_start_req, start_ack => Out_wrap_daemon_start_ack,  fin_req => Out_wrap_daemon_fin_req,  fin_ack => Out_wrap_daemon_fin_ack);
  -- module c_block_daemon
  c_block_daemon_instance:c_block_daemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => c_block_daemon_start_req,
      start_ack => c_block_daemon_start_ack,
      fin_req => c_block_daemon_fin_req,
      fin_ack => c_block_daemon_fin_ack,
      clk => clk,
      reset => reset,
      cmd_in_pipe_read_req => cmd_in_pipe_read_req(0 downto 0),
      cmd_in_pipe_read_ack => cmd_in_pipe_read_ack(0 downto 0),
      cmd_in_pipe_read_data => cmd_in_pipe_read_data(63 downto 0),
      d_block_done_pipe_read_req => d_block_done_pipe_read_req(0 downto 0),
      d_block_done_pipe_read_ack => d_block_done_pipe_read_ack(0 downto 0),
      d_block_done_pipe_read_data => d_block_done_pipe_read_data(0 downto 0),
      e_block_done_pipe_read_req => e_block_done_pipe_read_req(0 downto 0),
      e_block_done_pipe_read_ack => e_block_done_pipe_read_ack(0 downto 0),
      e_block_done_pipe_read_data => e_block_done_pipe_read_data(0 downto 0),
      d_cmd_pipe_pipe_write_req => d_cmd_pipe_pipe_write_req(0 downto 0),
      d_cmd_pipe_pipe_write_ack => d_cmd_pipe_pipe_write_ack(0 downto 0),
      d_cmd_pipe_pipe_write_data => d_cmd_pipe_pipe_write_data(143 downto 0),
      e_cmd_pipe_pipe_write_req => e_cmd_pipe_pipe_write_req(0 downto 0),
      e_cmd_pipe_pipe_write_ack => e_cmd_pipe_pipe_write_ack(0 downto 0),
      e_cmd_pipe_pipe_write_data => e_cmd_pipe_pipe_write_data(143 downto 0),
      status_out_pipe_write_req => status_out_pipe_write_req(0 downto 0),
      status_out_pipe_write_ack => status_out_pipe_write_ack(0 downto 0),
      status_out_pipe_write_data => status_out_pipe_write_data(63 downto 0),
      tag_in => c_block_daemon_tag_in,
      tag_out => c_block_daemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  c_block_daemon_tag_in <= (others => '0');
  c_block_daemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => c_block_daemon_start_req, start_ack => c_block_daemon_start_ack,  fin_req => c_block_daemon_fin_req,  fin_ack => c_block_daemon_fin_ack);
  -- module d_block_daemon
  d_block_daemon_instance:d_block_daemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => d_block_daemon_start_req,
      start_ack => d_block_daemon_start_ack,
      fin_req => d_block_daemon_fin_req,
      fin_ack => d_block_daemon_fin_ack,
      clk => clk,
      reset => reset,
      d_cmd_pipe_pipe_read_req => d_cmd_pipe_pipe_read_req(0 downto 0),
      d_cmd_pipe_pipe_read_ack => d_cmd_pipe_pipe_read_ack(0 downto 0),
      d_cmd_pipe_pipe_read_data => d_cmd_pipe_pipe_read_data(143 downto 0),
      d_in_buf_pipe_read_req => d_in_buf_pipe_read_req(0 downto 0),
      d_in_buf_pipe_read_ack => d_in_buf_pipe_read_ack(0 downto 0),
      d_in_buf_pipe_read_data => d_in_buf_pipe_read_data(127 downto 0),
      d_block_done_pipe_write_req => d_block_done_pipe_write_req(0 downto 0),
      d_block_done_pipe_write_ack => d_block_done_pipe_write_ack(0 downto 0),
      d_block_done_pipe_write_data => d_block_done_pipe_write_data(0 downto 0),
      d_out_buf_pipe_write_req => d_out_buf_pipe_write_req(0 downto 0),
      d_out_buf_pipe_write_ack => d_out_buf_pipe_write_ack(0 downto 0),
      d_out_buf_pipe_write_data => d_out_buf_pipe_write_data(127 downto 0),
      key_expand_single_call_reqs => key_expand_single_call_reqs(1 downto 1),
      key_expand_single_call_acks => key_expand_single_call_acks(1 downto 1),
      key_expand_single_call_data => key_expand_single_call_data(271 downto 136),
      key_expand_single_call_tag => key_expand_single_call_tag(7 downto 4),
      key_expand_single_return_reqs => key_expand_single_return_reqs(1 downto 1),
      key_expand_single_return_acks => key_expand_single_return_acks(1 downto 1),
      key_expand_single_return_data => key_expand_single_return_data(271 downto 136),
      key_expand_single_return_tag => key_expand_single_return_tag(7 downto 4),
      tag_in => d_block_daemon_tag_in,
      tag_out => d_block_daemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  d_block_daemon_tag_in <= (others => '0');
  d_block_daemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => d_block_daemon_start_req, start_ack => d_block_daemon_start_ack,  fin_req => d_block_daemon_fin_req,  fin_ack => d_block_daemon_fin_ack);
  -- module e_block_daemon
  e_block_daemon_instance:e_block_daemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => e_block_daemon_start_req,
      start_ack => e_block_daemon_start_ack,
      fin_req => e_block_daemon_fin_req,
      fin_ack => e_block_daemon_fin_ack,
      clk => clk,
      reset => reset,
      e_in_buf_pipe_read_req => e_in_buf_pipe_read_req(0 downto 0),
      e_in_buf_pipe_read_ack => e_in_buf_pipe_read_ack(0 downto 0),
      e_in_buf_pipe_read_data => e_in_buf_pipe_read_data(127 downto 0),
      e_cmd_pipe_pipe_read_req => e_cmd_pipe_pipe_read_req(0 downto 0),
      e_cmd_pipe_pipe_read_ack => e_cmd_pipe_pipe_read_ack(0 downto 0),
      e_cmd_pipe_pipe_read_data => e_cmd_pipe_pipe_read_data(143 downto 0),
      e_out_buf_pipe_write_req => e_out_buf_pipe_write_req(0 downto 0),
      e_out_buf_pipe_write_ack => e_out_buf_pipe_write_ack(0 downto 0),
      e_out_buf_pipe_write_data => e_out_buf_pipe_write_data(127 downto 0),
      e_block_done_pipe_write_req => e_block_done_pipe_write_req(0 downto 0),
      e_block_done_pipe_write_ack => e_block_done_pipe_write_ack(0 downto 0),
      e_block_done_pipe_write_data => e_block_done_pipe_write_data(0 downto 0),
      key_expand_single_call_reqs => key_expand_single_call_reqs(0 downto 0),
      key_expand_single_call_acks => key_expand_single_call_acks(0 downto 0),
      key_expand_single_call_data => key_expand_single_call_data(135 downto 0),
      key_expand_single_call_tag => key_expand_single_call_tag(3 downto 0),
      key_expand_single_return_reqs => key_expand_single_return_reqs(0 downto 0),
      key_expand_single_return_acks => key_expand_single_return_acks(0 downto 0),
      key_expand_single_return_data => key_expand_single_return_data(135 downto 0),
      key_expand_single_return_tag => key_expand_single_return_tag(3 downto 0),
      tag_in => e_block_daemon_tag_in,
      tag_out => e_block_daemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  e_block_daemon_tag_in <= (others => '0');
  e_block_daemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => e_block_daemon_start_req, start_ack => e_block_daemon_start_ack,  fin_req => e_block_daemon_fin_req,  fin_ack => e_block_daemon_fin_ack);
  -- module key_expand_single
  key_expand_single_K_in <= key_expand_single_in_args(135 downto 8);
  key_expand_single_Round_C <= key_expand_single_in_args(7 downto 0);
  key_expand_single_out_args <= key_expand_single_K_out & key_expand_single_nRound_C ;
  -- call arbiter for module key_expand_single
  key_expand_single_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 2,
      call_data_width => 136,
      return_data_width => 136,
      callee_tag_length => 2,
      caller_tag_length => 4--
    )
    port map(-- 
      call_reqs => key_expand_single_call_reqs,
      call_acks => key_expand_single_call_acks,
      return_reqs => key_expand_single_return_reqs,
      return_acks => key_expand_single_return_acks,
      call_data  => key_expand_single_call_data,
      call_tag  => key_expand_single_call_tag,
      return_tag  => key_expand_single_return_tag,
      call_mtag => key_expand_single_tag_in,
      return_mtag => key_expand_single_tag_out,
      return_data =>key_expand_single_return_data,
      call_mreq => key_expand_single_start_req,
      call_mack => key_expand_single_start_ack,
      return_mreq => key_expand_single_fin_req,
      return_mack => key_expand_single_fin_ack,
      call_mdata => key_expand_single_in_args,
      return_mdata => key_expand_single_out_args,
      clk => clk, 
      reset => reset --
    ); --
  key_expand_single_instance:key_expand_single-- 
    generic map(tag_length => 6)
    port map(-- 
      K_in => key_expand_single_K_in,
      Round_C => key_expand_single_Round_C,
      K_out => key_expand_single_K_out,
      nRound_C => key_expand_single_nRound_C,
      start_req => key_expand_single_start_req,
      start_ack => key_expand_single_start_ack,
      fin_req => key_expand_single_fin_req,
      fin_ack => key_expand_single_fin_ack,
      clk => clk,
      reset => reset,
      tag_in => key_expand_single_tag_in,
      tag_out => key_expand_single_tag_out-- 
    ); -- 
  -- module w_in_buff_daemon
  w_in_buff_daemon_instance:w_in_buff_daemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => w_in_buff_daemon_start_req,
      start_ack => w_in_buff_daemon_start_ack,
      fin_req => w_in_buff_daemon_fin_req,
      fin_ack => w_in_buff_daemon_fin_ack,
      clk => clk,
      reset => reset,
      in_data_pipe_read_req => in_data_pipe_read_req(0 downto 0),
      in_data_pipe_read_ack => in_data_pipe_read_ack(0 downto 0),
      in_data_pipe_read_data => in_data_pipe_read_data(63 downto 0),
      w_in_buf_pipe_write_req => w_in_buf_pipe_write_req(0 downto 0),
      w_in_buf_pipe_write_ack => w_in_buf_pipe_write_ack(0 downto 0),
      w_in_buf_pipe_write_data => w_in_buf_pipe_write_data(127 downto 0),
      tag_in => w_in_buff_daemon_tag_in,
      tag_out => w_in_buff_daemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  w_in_buff_daemon_tag_in <= (others => '0');
  w_in_buff_daemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => w_in_buff_daemon_start_req, start_ack => w_in_buff_daemon_start_ack,  fin_req => w_in_buff_daemon_fin_req,  fin_ack => w_in_buff_daemon_fin_ack);
  -- module w_out_buff_daemon
  w_out_buff_daemon_instance:w_out_buff_daemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => w_out_buff_daemon_start_req,
      start_ack => w_out_buff_daemon_start_ack,
      fin_req => w_out_buff_daemon_fin_req,
      fin_ack => w_out_buff_daemon_fin_ack,
      clk => clk,
      reset => reset,
      w_out_buf_pipe_read_req => w_out_buf_pipe_read_req(0 downto 0),
      w_out_buf_pipe_read_ack => w_out_buf_pipe_read_ack(0 downto 0),
      w_out_buf_pipe_read_data => w_out_buf_pipe_read_data(127 downto 0),
      out_data_pipe_write_req => out_data_pipe_write_req(0 downto 0),
      out_data_pipe_write_ack => out_data_pipe_write_ack(0 downto 0),
      out_data_pipe_write_data => out_data_pipe_write_data(63 downto 0),
      tag_in => w_out_buff_daemon_tag_in,
      tag_out => w_out_buff_daemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  w_out_buff_daemon_tag_in <= (others => '0');
  w_out_buff_daemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => w_out_buff_daemon_start_req, start_ack => w_out_buff_daemon_start_ack,  fin_req => w_out_buff_daemon_fin_req,  fin_ack => w_out_buff_daemon_fin_ack);
  cmd_in_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe cmd_in",
      num_reads => 1,
      num_writes => 1,
      data_width => 64,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      depth => 4 --
    )
    port map( -- 
      read_req => cmd_in_pipe_read_req,
      read_ack => cmd_in_pipe_read_ack,
      read_data => cmd_in_pipe_read_data,
      write_req => cmd_in_pipe_write_req,
      write_ack => cmd_in_pipe_write_ack,
      write_data => cmd_in_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  d_block_done_Pipe: NonBlockingReadPipeBase -- 
    generic map( -- 
      name => "pipe d_block_done",
      num_reads => 1,
      num_writes => 1,
      data_width => 1,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      depth => 2 --
    )
    port map( -- 
      read_req => d_block_done_pipe_read_req,
      read_ack => d_block_done_pipe_read_ack,
      read_data => d_block_done_pipe_read_data,
      write_req => d_block_done_pipe_write_req,
      write_ack => d_block_done_pipe_write_ack,
      write_data => d_block_done_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  d_cmd_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe d_cmd_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 144,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      depth => 2 --
    )
    port map( -- 
      read_req => d_cmd_pipe_pipe_read_req,
      read_ack => d_cmd_pipe_pipe_read_ack,
      read_data => d_cmd_pipe_pipe_read_data,
      write_req => d_cmd_pipe_pipe_write_req,
      write_ack => d_cmd_pipe_pipe_write_ack,
      write_data => d_cmd_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  d_in_buf_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe d_in_buf",
      num_reads => 1,
      num_writes => 1,
      data_width => 128,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      depth => 2 --
    )
    port map( -- 
      read_req => d_in_buf_pipe_read_req,
      read_ack => d_in_buf_pipe_read_ack,
      read_data => d_in_buf_pipe_read_data,
      write_req => d_in_buf_pipe_write_req,
      write_ack => d_in_buf_pipe_write_ack,
      write_data => d_in_buf_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  d_out_buf_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe d_out_buf",
      num_reads => 1,
      num_writes => 1,
      data_width => 128,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      depth => 2 --
    )
    port map( -- 
      read_req => d_out_buf_pipe_read_req,
      read_ack => d_out_buf_pipe_read_ack,
      read_data => d_out_buf_pipe_read_data,
      write_req => d_out_buf_pipe_write_req,
      write_ack => d_out_buf_pipe_write_ack,
      write_data => d_out_buf_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  e_block_done_Pipe: NonBlockingReadPipeBase -- 
    generic map( -- 
      name => "pipe e_block_done",
      num_reads => 1,
      num_writes => 1,
      data_width => 1,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      depth => 2 --
    )
    port map( -- 
      read_req => e_block_done_pipe_read_req,
      read_ack => e_block_done_pipe_read_ack,
      read_data => e_block_done_pipe_read_data,
      write_req => e_block_done_pipe_write_req,
      write_ack => e_block_done_pipe_write_ack,
      write_data => e_block_done_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  e_cmd_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe e_cmd_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 144,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      depth => 2 --
    )
    port map( -- 
      read_req => e_cmd_pipe_pipe_read_req,
      read_ack => e_cmd_pipe_pipe_read_ack,
      read_data => e_cmd_pipe_pipe_read_data,
      write_req => e_cmd_pipe_pipe_write_req,
      write_ack => e_cmd_pipe_pipe_write_ack,
      write_data => e_cmd_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  e_in_buf_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe e_in_buf",
      num_reads => 1,
      num_writes => 1,
      data_width => 128,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      depth => 2 --
    )
    port map( -- 
      read_req => e_in_buf_pipe_read_req,
      read_ack => e_in_buf_pipe_read_ack,
      read_data => e_in_buf_pipe_read_data,
      write_req => e_in_buf_pipe_write_req,
      write_ack => e_in_buf_pipe_write_ack,
      write_data => e_in_buf_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  e_out_buf_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe e_out_buf",
      num_reads => 1,
      num_writes => 1,
      data_width => 128,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      depth => 2 --
    )
    port map( -- 
      read_req => e_out_buf_pipe_read_req,
      read_ack => e_out_buf_pipe_read_ack,
      read_data => e_out_buf_pipe_read_data,
      write_req => e_out_buf_pipe_write_req,
      write_ack => e_out_buf_pipe_write_ack,
      write_data => e_out_buf_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  in_data_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe in_data",
      num_reads => 1,
      num_writes => 1,
      data_width => 64,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      depth => 2 --
    )
    port map( -- 
      read_req => in_data_pipe_read_req,
      read_ack => in_data_pipe_read_ack,
      read_data => in_data_pipe_read_data,
      write_req => in_data_pipe_write_req,
      write_ack => in_data_pipe_write_ack,
      write_data => in_data_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  out_data_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe out_data",
      num_reads => 1,
      num_writes => 1,
      data_width => 64,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      depth => 2 --
    )
    port map( -- 
      read_req => out_data_pipe_read_req,
      read_ack => out_data_pipe_read_ack,
      read_data => out_data_pipe_read_data,
      write_req => out_data_pipe_write_req,
      write_ack => out_data_pipe_write_ack,
      write_data => out_data_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  out_wrap_cmd_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe out_wrap_cmd",
      num_reads => 1,
      num_writes => 1,
      data_width => 64,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      depth => 2 --
    )
    port map( -- 
      read_req => out_wrap_cmd_pipe_read_req,
      read_ack => out_wrap_cmd_pipe_read_ack,
      read_data => out_wrap_cmd_pipe_read_data,
      write_req => out_wrap_cmd_pipe_write_req,
      write_ack => out_wrap_cmd_pipe_write_ack,
      write_data => out_wrap_cmd_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  out_wrap_data_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe out_wrap_data",
      num_reads => 1,
      num_writes => 1,
      data_width => 128,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      depth => 2 --
    )
    port map( -- 
      read_req => out_wrap_data_pipe_read_req,
      read_ack => out_wrap_data_pipe_read_ack,
      read_data => out_wrap_data_pipe_read_data,
      write_req => out_wrap_data_pipe_write_req,
      write_ack => out_wrap_data_pipe_write_ack,
      write_data => out_wrap_data_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  status_out_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe status_out",
      num_reads => 1,
      num_writes => 1,
      data_width => 64,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      depth => 2 --
    )
    port map( -- 
      read_req => status_out_pipe_read_req,
      read_ack => status_out_pipe_read_ack,
      read_data => status_out_pipe_read_data,
      write_req => status_out_pipe_write_req,
      write_ack => status_out_pipe_write_ack,
      write_data => status_out_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  w_in_buf_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe w_in_buf",
      num_reads => 1,
      num_writes => 1,
      data_width => 128,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      depth => 512 --
    )
    port map( -- 
      read_req => w_in_buf_pipe_read_req,
      read_ack => w_in_buf_pipe_read_ack,
      read_data => w_in_buf_pipe_read_data,
      write_req => w_in_buf_pipe_write_req,
      write_ack => w_in_buf_pipe_write_ack,
      write_data => w_in_buf_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  w_out_buf_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe w_out_buf",
      num_reads => 1,
      num_writes => 1,
      data_width => 128,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      depth => 512 --
    )
    port map( -- 
      read_req => w_out_buf_pipe_read_req,
      read_ack => w_out_buf_pipe_read_ack,
      read_data => w_out_buf_pipe_read_data,
      write_req => w_out_buf_pipe_write_req,
      write_ack => w_out_buf_pipe_write_ack,
      write_data => w_out_buf_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- 
end ahir_system_arch;
